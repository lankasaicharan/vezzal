magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 654 241 1136 263
rect 56 49 1136 241
rect 0 0 1152 49
<< scnmos >>
rect 135 47 165 215
rect 221 47 251 215
rect 307 47 337 215
rect 393 47 423 215
rect 479 47 509 215
rect 737 69 767 237
rect 823 69 853 237
rect 925 69 955 237
rect 1027 69 1057 237
<< scpmoshvt >>
rect 97 367 127 619
rect 221 367 251 619
rect 307 367 337 619
rect 425 367 455 619
rect 511 367 541 619
rect 737 367 767 619
rect 823 367 853 619
rect 909 367 939 619
rect 995 367 1025 619
<< ndiff >>
rect 680 229 737 237
rect 82 203 135 215
rect 82 169 90 203
rect 124 169 135 203
rect 82 101 135 169
rect 82 67 90 101
rect 124 67 135 101
rect 82 47 135 67
rect 165 163 221 215
rect 165 129 176 163
rect 210 129 221 163
rect 165 89 221 129
rect 165 55 176 89
rect 210 55 221 89
rect 165 47 221 55
rect 251 203 307 215
rect 251 169 262 203
rect 296 169 307 203
rect 251 101 307 169
rect 251 67 262 101
rect 296 67 307 101
rect 251 47 307 67
rect 337 161 393 215
rect 337 127 348 161
rect 382 127 393 161
rect 337 93 393 127
rect 337 59 348 93
rect 382 59 393 93
rect 337 47 393 59
rect 423 93 479 215
rect 423 59 434 93
rect 468 59 479 93
rect 423 47 479 59
rect 509 173 562 215
rect 509 139 520 173
rect 554 139 562 173
rect 509 47 562 139
rect 680 195 692 229
rect 726 195 737 229
rect 680 69 737 195
rect 767 159 823 237
rect 767 125 778 159
rect 812 125 823 159
rect 767 69 823 125
rect 853 225 925 237
rect 853 191 880 225
rect 914 191 925 225
rect 853 155 925 191
rect 853 121 880 155
rect 914 121 925 155
rect 853 69 925 121
rect 955 181 1027 237
rect 955 147 982 181
rect 1016 147 1027 181
rect 955 111 1027 147
rect 955 77 982 111
rect 1016 77 1027 111
rect 955 69 1027 77
rect 1057 225 1110 237
rect 1057 191 1068 225
rect 1102 191 1110 225
rect 1057 116 1110 191
rect 1057 82 1068 116
rect 1102 82 1110 116
rect 1057 69 1110 82
<< pdiff >>
rect 352 626 410 638
rect 352 619 364 626
rect 44 599 97 619
rect 44 565 52 599
rect 86 565 97 599
rect 44 504 97 565
rect 44 470 52 504
rect 86 470 97 504
rect 44 413 97 470
rect 44 379 52 413
rect 86 379 97 413
rect 44 367 97 379
rect 127 607 221 619
rect 127 573 158 607
rect 192 573 221 607
rect 127 492 221 573
rect 127 458 158 492
rect 192 458 221 492
rect 127 367 221 458
rect 251 594 307 619
rect 251 560 262 594
rect 296 560 307 594
rect 251 492 307 560
rect 251 458 262 492
rect 296 458 307 492
rect 251 367 307 458
rect 337 592 364 619
rect 398 619 410 626
rect 563 626 621 638
rect 563 619 575 626
rect 398 592 425 619
rect 337 367 425 592
rect 455 486 511 619
rect 455 452 466 486
rect 500 452 511 486
rect 455 418 511 452
rect 455 384 466 418
rect 500 384 511 418
rect 455 367 511 384
rect 541 592 575 619
rect 609 592 621 626
rect 541 367 621 592
rect 684 416 737 619
rect 684 382 692 416
rect 726 382 737 416
rect 684 367 737 382
rect 767 531 823 619
rect 767 497 778 531
rect 812 497 823 531
rect 767 367 823 497
rect 853 544 909 619
rect 853 510 864 544
rect 898 510 909 544
rect 853 436 909 510
rect 853 402 864 436
rect 898 402 909 436
rect 853 367 909 402
rect 939 599 995 619
rect 939 565 950 599
rect 984 565 995 599
rect 939 504 995 565
rect 939 470 950 504
rect 984 470 995 504
rect 939 367 995 470
rect 1025 599 1078 619
rect 1025 565 1036 599
rect 1070 565 1078 599
rect 1025 509 1078 565
rect 1025 475 1036 509
rect 1070 475 1078 509
rect 1025 418 1078 475
rect 1025 384 1036 418
rect 1070 384 1078 418
rect 1025 367 1078 384
<< ndiffc >>
rect 90 169 124 203
rect 90 67 124 101
rect 176 129 210 163
rect 176 55 210 89
rect 262 169 296 203
rect 262 67 296 101
rect 348 127 382 161
rect 348 59 382 93
rect 434 59 468 93
rect 520 139 554 173
rect 692 195 726 229
rect 778 125 812 159
rect 880 191 914 225
rect 880 121 914 155
rect 982 147 1016 181
rect 982 77 1016 111
rect 1068 191 1102 225
rect 1068 82 1102 116
<< pdiffc >>
rect 52 565 86 599
rect 52 470 86 504
rect 52 379 86 413
rect 158 573 192 607
rect 158 458 192 492
rect 262 560 296 594
rect 262 458 296 492
rect 364 592 398 626
rect 466 452 500 486
rect 466 384 500 418
rect 575 592 609 626
rect 692 382 726 416
rect 778 497 812 531
rect 864 510 898 544
rect 864 402 898 436
rect 950 565 984 599
rect 950 470 984 504
rect 1036 565 1070 599
rect 1036 475 1070 509
rect 1036 384 1070 418
<< poly >>
rect 97 619 127 645
rect 221 619 251 645
rect 307 619 337 645
rect 425 619 455 645
rect 511 619 541 645
rect 737 619 767 645
rect 823 619 853 645
rect 909 619 939 645
rect 995 619 1025 645
rect 97 335 127 367
rect 97 319 172 335
rect 97 285 122 319
rect 156 285 172 319
rect 97 269 172 285
rect 221 333 251 367
rect 307 333 337 367
rect 425 335 455 367
rect 221 317 337 333
rect 221 283 237 317
rect 271 283 337 317
rect 135 215 165 269
rect 221 267 337 283
rect 389 319 455 335
rect 389 285 405 319
rect 439 299 455 319
rect 511 299 541 367
rect 439 285 541 299
rect 389 269 541 285
rect 737 335 767 367
rect 823 335 853 367
rect 737 319 853 335
rect 737 285 803 319
rect 837 285 853 319
rect 737 269 853 285
rect 909 299 939 367
rect 995 335 1025 367
rect 991 319 1057 335
rect 991 299 1007 319
rect 909 285 1007 299
rect 1041 285 1057 319
rect 909 269 1057 285
rect 221 215 251 267
rect 307 215 337 267
rect 393 215 423 269
rect 479 215 509 269
rect 737 237 767 269
rect 823 237 853 269
rect 925 237 955 269
rect 1027 237 1057 269
rect 135 21 165 47
rect 221 21 251 47
rect 307 21 337 47
rect 393 21 423 47
rect 479 21 509 47
rect 737 43 767 69
rect 823 43 853 69
rect 925 43 955 69
rect 1027 43 1057 69
<< polycont >>
rect 122 285 156 319
rect 237 283 271 317
rect 405 285 439 319
rect 803 285 837 319
rect 1007 285 1041 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 36 599 88 615
rect 36 565 52 599
rect 86 565 88 599
rect 36 504 88 565
rect 36 470 52 504
rect 86 470 88 504
rect 36 413 88 470
rect 142 607 208 649
rect 142 573 158 607
rect 192 573 208 607
rect 348 626 414 649
rect 142 492 208 573
rect 142 458 158 492
rect 192 458 208 492
rect 246 560 262 594
rect 296 560 312 594
rect 348 592 364 626
rect 398 592 414 626
rect 348 588 414 592
rect 559 626 625 649
rect 559 592 575 626
rect 609 592 625 626
rect 559 588 625 592
rect 661 599 993 615
rect 246 554 312 560
rect 661 581 950 599
rect 661 554 695 581
rect 246 520 695 554
rect 948 565 950 581
rect 984 565 993 599
rect 762 531 814 547
rect 246 492 312 520
rect 246 458 262 492
rect 296 458 312 492
rect 762 497 778 531
rect 812 497 814 531
rect 762 486 814 497
rect 450 452 466 486
rect 500 452 814 486
rect 848 544 914 547
rect 848 510 864 544
rect 898 510 914 544
rect 36 379 52 413
rect 86 379 88 413
rect 36 231 88 379
rect 122 371 370 424
rect 122 319 158 371
rect 156 285 158 319
rect 336 334 370 371
rect 450 418 516 452
rect 848 436 914 510
rect 948 504 993 565
rect 948 470 950 504
rect 984 470 993 504
rect 948 454 993 470
rect 1027 599 1086 615
rect 1027 565 1036 599
rect 1070 565 1086 599
rect 1027 509 1086 565
rect 1027 475 1036 509
rect 1070 475 1086 509
rect 848 418 864 436
rect 450 384 466 418
rect 500 384 516 418
rect 450 368 516 384
rect 574 416 864 418
rect 574 382 692 416
rect 726 402 864 416
rect 898 420 914 436
rect 1027 420 1086 475
rect 898 418 1086 420
rect 898 402 1036 418
rect 726 384 1036 402
rect 1070 384 1086 418
rect 726 382 742 384
rect 336 319 455 334
rect 122 269 158 285
rect 192 283 237 317
rect 271 283 287 317
rect 336 285 405 319
rect 439 285 455 319
rect 574 316 742 382
rect 192 231 226 283
rect 336 281 455 285
rect 676 249 742 316
rect 787 319 943 350
rect 787 285 803 319
rect 837 285 943 319
rect 977 319 1134 350
rect 977 285 1007 319
rect 1041 285 1134 319
rect 36 203 226 231
rect 36 169 90 203
rect 124 197 226 203
rect 260 213 642 247
rect 260 203 306 213
rect 124 169 126 197
rect 36 101 126 169
rect 260 169 262 203
rect 296 169 306 203
rect 36 67 90 101
rect 124 67 126 101
rect 36 51 126 67
rect 160 129 176 163
rect 210 129 226 163
rect 160 89 226 129
rect 160 55 176 89
rect 210 55 226 89
rect 160 17 226 55
rect 260 101 306 169
rect 260 67 262 101
rect 296 67 306 101
rect 260 51 306 67
rect 340 173 570 179
rect 340 161 520 173
rect 340 127 348 161
rect 382 139 520 161
rect 554 139 570 173
rect 382 135 570 139
rect 604 159 642 213
rect 676 229 1118 249
rect 676 195 692 229
rect 726 225 1118 229
rect 726 195 880 225
rect 676 193 880 195
rect 864 191 880 193
rect 914 215 1068 225
rect 914 191 930 215
rect 382 127 384 135
rect 340 93 384 127
rect 604 125 778 159
rect 812 125 828 159
rect 604 121 828 125
rect 864 155 930 191
rect 1066 191 1068 215
rect 1102 191 1118 225
rect 864 121 880 155
rect 914 121 930 155
rect 966 147 982 181
rect 1016 147 1032 181
rect 966 111 1032 147
rect 340 59 348 93
rect 382 59 384 93
rect 340 17 384 59
rect 418 93 484 101
rect 418 59 434 93
rect 468 87 484 93
rect 966 87 982 111
rect 468 77 982 87
rect 1016 77 1032 111
rect 468 59 1032 77
rect 1066 116 1118 191
rect 1066 82 1068 116
rect 1102 82 1118 116
rect 1066 66 1118 82
rect 418 51 1032 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3849140
string GDS_START 3840040
<< end >>
