magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 17 243 957 259
rect 17 49 1235 243
rect 0 0 1248 49
<< scnmos >>
rect 96 65 126 233
rect 182 65 212 233
rect 268 65 298 233
rect 354 65 384 233
rect 576 65 606 233
rect 662 65 692 233
rect 748 65 778 233
rect 834 65 864 233
rect 1040 49 1070 217
rect 1126 49 1156 217
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 268 367 298 619
rect 354 367 384 619
rect 487 367 517 619
rect 662 367 692 619
rect 764 367 794 619
rect 924 367 954 619
rect 1010 367 1040 619
rect 1096 367 1126 619
<< ndiff >>
rect 43 192 96 233
rect 43 158 51 192
rect 85 158 96 192
rect 43 113 96 158
rect 43 79 51 113
rect 85 79 96 113
rect 43 65 96 79
rect 126 132 182 233
rect 126 98 137 132
rect 171 98 182 132
rect 126 65 182 98
rect 212 192 268 233
rect 212 158 223 192
rect 257 158 268 192
rect 212 111 268 158
rect 212 77 223 111
rect 257 77 268 111
rect 212 65 268 77
rect 298 225 354 233
rect 298 191 309 225
rect 343 191 354 225
rect 298 155 354 191
rect 298 121 309 155
rect 343 121 354 155
rect 298 65 354 121
rect 384 181 451 233
rect 384 147 409 181
rect 443 147 451 181
rect 384 111 451 147
rect 384 77 409 111
rect 443 77 451 111
rect 384 65 451 77
rect 509 181 576 233
rect 509 147 517 181
rect 551 147 576 181
rect 509 111 576 147
rect 509 77 517 111
rect 551 77 576 111
rect 509 65 576 77
rect 606 225 662 233
rect 606 191 617 225
rect 651 191 662 225
rect 606 155 662 191
rect 606 121 617 155
rect 651 121 662 155
rect 606 65 662 121
rect 692 225 748 233
rect 692 191 703 225
rect 737 191 748 225
rect 692 111 748 191
rect 692 77 703 111
rect 737 77 748 111
rect 692 65 748 77
rect 778 225 834 233
rect 778 191 789 225
rect 823 191 834 225
rect 778 155 834 191
rect 778 121 789 155
rect 823 121 834 155
rect 778 65 834 121
rect 864 181 931 233
rect 864 147 889 181
rect 923 147 931 181
rect 864 111 931 147
rect 864 77 889 111
rect 923 77 931 111
rect 864 65 931 77
rect 987 181 1040 217
rect 987 147 995 181
rect 1029 147 1040 181
rect 987 95 1040 147
rect 987 61 995 95
rect 1029 61 1040 95
rect 987 49 1040 61
rect 1070 205 1126 217
rect 1070 171 1081 205
rect 1115 171 1126 205
rect 1070 101 1126 171
rect 1070 67 1081 101
rect 1115 67 1126 101
rect 1070 49 1126 67
rect 1156 205 1209 217
rect 1156 171 1167 205
rect 1201 171 1209 205
rect 1156 95 1209 171
rect 1156 61 1167 95
rect 1201 61 1209 95
rect 1156 49 1209 61
<< pdiff >>
rect 43 599 96 619
rect 43 565 51 599
rect 85 565 96 599
rect 43 515 96 565
rect 43 481 51 515
rect 85 481 96 515
rect 43 436 96 481
rect 43 402 51 436
rect 85 402 96 436
rect 43 367 96 402
rect 126 547 182 619
rect 126 513 137 547
rect 171 513 182 547
rect 126 479 182 513
rect 126 445 137 479
rect 171 445 182 479
rect 126 411 182 445
rect 126 377 137 411
rect 171 377 182 411
rect 126 367 182 377
rect 212 597 268 619
rect 212 563 223 597
rect 257 563 268 597
rect 212 529 268 563
rect 212 495 223 529
rect 257 495 268 529
rect 212 457 268 495
rect 212 423 223 457
rect 257 423 268 457
rect 212 367 268 423
rect 298 547 354 619
rect 298 513 309 547
rect 343 513 354 547
rect 298 479 354 513
rect 298 445 309 479
rect 343 445 354 479
rect 298 411 354 445
rect 298 377 309 411
rect 343 377 354 411
rect 298 367 354 377
rect 384 608 487 619
rect 384 574 419 608
rect 453 574 487 608
rect 384 498 487 574
rect 384 464 419 498
rect 453 464 487 498
rect 384 367 487 464
rect 517 569 662 619
rect 517 535 528 569
rect 562 535 617 569
rect 651 535 662 569
rect 517 367 662 535
rect 692 599 764 619
rect 692 565 711 599
rect 745 565 764 599
rect 692 514 764 565
rect 692 480 711 514
rect 745 480 764 514
rect 692 434 764 480
rect 692 400 711 434
rect 745 400 764 434
rect 692 367 764 400
rect 794 607 924 619
rect 794 573 805 607
rect 839 573 879 607
rect 913 573 924 607
rect 794 494 924 573
rect 794 460 805 494
rect 839 460 879 494
rect 913 460 924 494
rect 794 367 924 460
rect 954 599 1010 619
rect 954 565 965 599
rect 999 565 1010 599
rect 954 506 1010 565
rect 954 472 965 506
rect 999 472 1010 506
rect 954 413 1010 472
rect 954 379 965 413
rect 999 379 1010 413
rect 954 367 1010 379
rect 1040 607 1096 619
rect 1040 573 1051 607
rect 1085 573 1096 607
rect 1040 531 1096 573
rect 1040 497 1051 531
rect 1085 497 1096 531
rect 1040 453 1096 497
rect 1040 419 1051 453
rect 1085 419 1096 453
rect 1040 367 1096 419
rect 1126 599 1179 619
rect 1126 565 1137 599
rect 1171 565 1179 599
rect 1126 503 1179 565
rect 1126 469 1137 503
rect 1171 469 1179 503
rect 1126 413 1179 469
rect 1126 379 1137 413
rect 1171 379 1179 413
rect 1126 367 1179 379
<< ndiffc >>
rect 51 158 85 192
rect 51 79 85 113
rect 137 98 171 132
rect 223 158 257 192
rect 223 77 257 111
rect 309 191 343 225
rect 309 121 343 155
rect 409 147 443 181
rect 409 77 443 111
rect 517 147 551 181
rect 517 77 551 111
rect 617 191 651 225
rect 617 121 651 155
rect 703 191 737 225
rect 703 77 737 111
rect 789 191 823 225
rect 789 121 823 155
rect 889 147 923 181
rect 889 77 923 111
rect 995 147 1029 181
rect 995 61 1029 95
rect 1081 171 1115 205
rect 1081 67 1115 101
rect 1167 171 1201 205
rect 1167 61 1201 95
<< pdiffc >>
rect 51 565 85 599
rect 51 481 85 515
rect 51 402 85 436
rect 137 513 171 547
rect 137 445 171 479
rect 137 377 171 411
rect 223 563 257 597
rect 223 495 257 529
rect 223 423 257 457
rect 309 513 343 547
rect 309 445 343 479
rect 309 377 343 411
rect 419 574 453 608
rect 419 464 453 498
rect 528 535 562 569
rect 617 535 651 569
rect 711 565 745 599
rect 711 480 745 514
rect 711 400 745 434
rect 805 573 839 607
rect 879 573 913 607
rect 805 460 839 494
rect 879 460 913 494
rect 965 565 999 599
rect 965 472 999 506
rect 965 379 999 413
rect 1051 573 1085 607
rect 1051 497 1085 531
rect 1051 419 1085 453
rect 1137 565 1171 599
rect 1137 469 1171 503
rect 1137 379 1171 413
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 268 619 298 645
rect 354 619 384 645
rect 487 619 517 645
rect 662 619 692 645
rect 764 619 794 645
rect 924 619 954 645
rect 1010 619 1040 645
rect 1096 619 1126 645
rect 96 321 126 367
rect 182 321 212 367
rect 47 305 212 321
rect 47 271 63 305
rect 97 271 162 305
rect 196 271 212 305
rect 47 255 212 271
rect 96 233 126 255
rect 182 233 212 255
rect 268 299 298 367
rect 354 335 384 367
rect 487 335 517 367
rect 662 335 692 367
rect 764 335 794 367
rect 924 335 954 367
rect 354 319 445 335
rect 354 299 395 319
rect 268 285 395 299
rect 429 285 445 319
rect 268 269 445 285
rect 487 319 692 335
rect 487 285 503 319
rect 537 285 692 319
rect 487 269 692 285
rect 268 233 298 269
rect 354 233 384 269
rect 576 233 606 269
rect 662 233 692 269
rect 748 319 954 335
rect 748 285 764 319
rect 798 285 881 319
rect 915 285 954 319
rect 748 269 954 285
rect 1010 305 1040 367
rect 1096 305 1126 367
rect 1010 289 1201 305
rect 748 233 778 269
rect 834 233 864 269
rect 1010 255 1151 289
rect 1185 255 1201 289
rect 1010 239 1201 255
rect 1040 217 1070 239
rect 1126 217 1156 239
rect 96 39 126 65
rect 182 39 212 65
rect 268 39 298 65
rect 354 39 384 65
rect 576 39 606 65
rect 662 39 692 65
rect 748 39 778 65
rect 834 39 864 65
rect 1040 23 1070 49
rect 1126 23 1156 49
<< polycont >>
rect 63 271 97 305
rect 162 271 196 305
rect 395 285 429 319
rect 503 285 537 319
rect 764 285 798 319
rect 881 285 915 319
rect 1151 255 1185 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 35 608 469 615
rect 35 599 419 608
rect 35 565 51 599
rect 85 597 419 599
rect 85 581 223 597
rect 85 565 87 581
rect 35 515 87 565
rect 221 563 223 581
rect 257 581 419 597
rect 257 563 259 581
rect 35 481 51 515
rect 85 481 87 515
rect 35 436 87 481
rect 35 402 51 436
rect 85 402 87 436
rect 35 386 87 402
rect 121 513 137 547
rect 171 513 187 547
rect 121 479 187 513
rect 121 445 137 479
rect 171 445 187 479
rect 121 411 187 445
rect 121 377 137 411
rect 171 377 187 411
rect 221 529 259 563
rect 403 574 419 581
rect 453 574 469 608
rect 221 495 223 529
rect 257 495 259 529
rect 221 457 259 495
rect 221 423 223 457
rect 257 423 259 457
rect 221 407 259 423
rect 293 513 309 547
rect 343 513 359 547
rect 293 479 359 513
rect 293 445 309 479
rect 343 445 359 479
rect 403 498 469 574
rect 512 569 667 649
rect 512 535 528 569
rect 562 535 617 569
rect 651 535 667 569
rect 512 526 667 535
rect 701 599 755 615
rect 701 565 711 599
rect 745 565 755 599
rect 403 464 419 498
rect 453 492 469 498
rect 701 514 755 565
rect 701 492 711 514
rect 453 480 711 492
rect 745 480 755 514
rect 453 464 755 480
rect 403 458 755 464
rect 293 424 359 445
rect 703 434 755 458
rect 789 607 929 649
rect 789 573 805 607
rect 839 573 879 607
rect 913 573 929 607
rect 789 494 929 573
rect 789 460 805 494
rect 839 460 879 494
rect 913 460 929 494
rect 789 452 929 460
rect 963 599 1001 615
rect 963 565 965 599
rect 999 565 1001 599
rect 963 506 1001 565
rect 963 472 965 506
rect 999 472 1001 506
rect 293 411 667 424
rect 121 373 187 377
rect 293 377 309 411
rect 343 384 667 411
rect 703 400 711 434
rect 745 418 755 434
rect 963 418 1001 472
rect 1035 607 1101 649
rect 1035 573 1051 607
rect 1085 573 1101 607
rect 1035 531 1101 573
rect 1035 497 1051 531
rect 1085 497 1101 531
rect 1035 453 1101 497
rect 1035 419 1051 453
rect 1085 419 1101 453
rect 1135 599 1187 615
rect 1135 565 1137 599
rect 1171 565 1187 599
rect 1135 503 1187 565
rect 1135 469 1137 503
rect 1171 469 1187 503
rect 745 413 1001 418
rect 745 400 965 413
rect 703 384 965 400
rect 343 377 345 384
rect 293 373 345 377
rect 17 305 87 352
rect 121 339 345 373
rect 379 319 453 350
rect 17 271 63 305
rect 97 271 162 305
rect 196 271 212 305
rect 379 285 395 319
rect 429 285 453 319
rect 487 319 553 350
rect 487 285 503 319
rect 537 285 553 319
rect 17 255 212 271
rect 17 242 97 255
rect 601 249 667 384
rect 999 385 1001 413
rect 1135 413 1187 469
rect 1135 385 1137 413
rect 999 379 1137 385
rect 1171 379 1187 413
rect 965 351 1187 379
rect 703 319 931 350
rect 703 285 764 319
rect 798 285 881 319
rect 915 285 931 319
rect 1151 289 1231 305
rect 1185 255 1231 289
rect 293 225 667 249
rect 35 192 259 208
rect 35 158 51 192
rect 85 174 223 192
rect 85 158 87 174
rect 35 113 87 158
rect 221 158 223 174
rect 257 158 259 192
rect 35 79 51 113
rect 85 79 87 113
rect 35 63 87 79
rect 121 132 187 140
rect 121 98 137 132
rect 171 98 187 132
rect 121 17 187 98
rect 221 111 259 158
rect 293 191 309 225
rect 343 215 617 225
rect 343 191 359 215
rect 293 155 359 191
rect 601 191 617 215
rect 651 191 667 225
rect 293 121 309 155
rect 343 121 359 155
rect 393 147 409 181
rect 443 147 459 181
rect 221 77 223 111
rect 257 87 259 111
rect 393 111 459 147
rect 393 87 409 111
rect 257 77 409 87
rect 443 77 459 111
rect 221 53 459 77
rect 501 147 517 181
rect 551 147 567 181
rect 501 111 567 147
rect 601 155 667 191
rect 601 121 617 155
rect 651 121 667 155
rect 701 225 739 241
rect 701 191 703 225
rect 737 191 739 225
rect 501 77 517 111
rect 551 87 567 111
rect 701 111 739 191
rect 773 225 1117 249
rect 1151 239 1231 255
rect 773 191 789 225
rect 823 215 1117 225
rect 823 191 839 215
rect 773 155 839 191
rect 1079 205 1117 215
rect 773 121 789 155
rect 823 121 839 155
rect 873 147 889 181
rect 923 147 939 181
rect 701 87 703 111
rect 551 77 703 87
rect 737 87 739 111
rect 873 111 939 147
rect 873 87 889 111
rect 737 77 889 87
rect 923 77 939 111
rect 501 53 939 77
rect 979 147 995 181
rect 1029 147 1045 181
rect 979 95 1045 147
rect 979 61 995 95
rect 1029 61 1045 95
rect 979 17 1045 61
rect 1079 171 1081 205
rect 1115 171 1117 205
rect 1079 101 1117 171
rect 1079 67 1081 101
rect 1115 67 1117 101
rect 1079 51 1117 67
rect 1151 171 1167 205
rect 1201 171 1217 205
rect 1151 95 1217 171
rect 1151 61 1167 95
rect 1201 61 1217 95
rect 1151 17 1217 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32oi_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1038588
string GDS_START 1027526
<< end >>
