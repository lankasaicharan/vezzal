magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 1 242 1418 248
rect 1 49 1439 242
rect 0 0 1440 49
<< scpmos >>
rect 86 368 116 536
rect 191 368 221 592
rect 393 368 423 592
rect 483 368 513 592
rect 573 368 603 592
rect 673 368 703 592
rect 773 368 803 592
rect 863 368 893 592
rect 953 368 983 592
rect 1044 368 1074 592
rect 1134 368 1164 592
rect 1224 368 1254 592
rect 1314 368 1344 592
<< nmoslvt >>
rect 84 112 114 222
rect 200 74 230 222
rect 398 74 428 222
rect 484 74 514 222
rect 570 74 600 222
rect 670 74 700 222
rect 756 74 786 222
rect 856 74 886 222
rect 942 74 972 222
rect 1028 74 1058 222
rect 1126 74 1156 222
rect 1226 74 1256 222
rect 1312 74 1342 222
<< ndiff >>
rect 27 184 84 222
rect 27 150 39 184
rect 73 150 84 184
rect 27 112 84 150
rect 114 152 200 222
rect 114 118 141 152
rect 175 118 200 152
rect 114 112 200 118
rect 129 74 200 112
rect 230 210 287 222
rect 230 176 241 210
rect 275 176 287 210
rect 230 120 287 176
rect 230 86 241 120
rect 275 86 287 120
rect 230 74 287 86
rect 341 210 398 222
rect 341 176 353 210
rect 387 176 398 210
rect 341 120 398 176
rect 341 86 353 120
rect 387 86 398 120
rect 341 74 398 86
rect 428 126 484 222
rect 428 92 439 126
rect 473 92 484 126
rect 428 74 484 92
rect 514 210 570 222
rect 514 176 525 210
rect 559 176 570 210
rect 514 74 570 176
rect 600 126 670 222
rect 600 92 611 126
rect 645 92 670 126
rect 600 74 670 92
rect 700 210 756 222
rect 700 176 711 210
rect 745 176 756 210
rect 700 120 756 176
rect 700 86 711 120
rect 745 86 756 120
rect 700 74 756 86
rect 786 126 856 222
rect 786 92 811 126
rect 845 92 856 126
rect 786 74 856 92
rect 886 210 942 222
rect 886 176 897 210
rect 931 176 942 210
rect 886 74 942 176
rect 972 126 1028 222
rect 972 92 983 126
rect 1017 92 1028 126
rect 972 74 1028 92
rect 1058 210 1126 222
rect 1058 176 1075 210
rect 1109 176 1126 210
rect 1058 74 1126 176
rect 1156 126 1226 222
rect 1156 92 1167 126
rect 1201 92 1226 126
rect 1156 74 1226 92
rect 1256 210 1312 222
rect 1256 176 1267 210
rect 1301 176 1312 210
rect 1256 120 1312 176
rect 1256 86 1267 120
rect 1301 86 1312 120
rect 1256 74 1312 86
rect 1342 216 1392 222
rect 1342 204 1413 216
rect 1342 170 1367 204
rect 1401 170 1413 204
rect 1342 120 1413 170
rect 1342 86 1367 120
rect 1401 86 1413 120
rect 1342 74 1413 86
<< pdiff >>
rect 138 536 191 592
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 429 86 490
rect 27 395 39 429
rect 73 395 86 429
rect 27 368 86 395
rect 116 524 191 536
rect 116 490 131 524
rect 165 490 191 524
rect 116 368 191 490
rect 221 580 280 592
rect 221 546 234 580
rect 268 546 280 580
rect 221 497 280 546
rect 221 463 234 497
rect 268 463 280 497
rect 221 414 280 463
rect 221 380 234 414
rect 268 380 280 414
rect 221 368 280 380
rect 334 580 393 592
rect 334 546 346 580
rect 380 546 393 580
rect 334 497 393 546
rect 334 463 346 497
rect 380 463 393 497
rect 334 414 393 463
rect 334 380 346 414
rect 380 380 393 414
rect 334 368 393 380
rect 423 580 483 592
rect 423 546 436 580
rect 470 546 483 580
rect 423 482 483 546
rect 423 448 436 482
rect 470 448 483 482
rect 423 368 483 448
rect 513 580 573 592
rect 513 546 526 580
rect 560 546 573 580
rect 513 497 573 546
rect 513 463 526 497
rect 560 463 573 497
rect 513 414 573 463
rect 513 380 526 414
rect 560 380 573 414
rect 513 368 573 380
rect 603 580 673 592
rect 603 546 626 580
rect 660 546 673 580
rect 603 497 673 546
rect 603 463 626 497
rect 660 463 673 497
rect 603 414 673 463
rect 603 380 626 414
rect 660 380 673 414
rect 603 368 673 380
rect 703 580 773 592
rect 703 546 726 580
rect 760 546 773 580
rect 703 497 773 546
rect 703 463 726 497
rect 760 463 773 497
rect 703 414 773 463
rect 703 380 726 414
rect 760 380 773 414
rect 703 368 773 380
rect 803 580 863 592
rect 803 546 816 580
rect 850 546 863 580
rect 803 478 863 546
rect 803 444 816 478
rect 850 444 863 478
rect 803 368 863 444
rect 893 580 953 592
rect 893 546 906 580
rect 940 546 953 580
rect 893 497 953 546
rect 893 463 906 497
rect 940 463 953 497
rect 893 414 953 463
rect 893 380 906 414
rect 940 380 953 414
rect 893 368 953 380
rect 983 580 1044 592
rect 983 546 996 580
rect 1030 546 1044 580
rect 983 478 1044 546
rect 983 444 996 478
rect 1030 444 1044 478
rect 983 368 1044 444
rect 1074 580 1134 592
rect 1074 546 1087 580
rect 1121 546 1134 580
rect 1074 497 1134 546
rect 1074 463 1087 497
rect 1121 463 1134 497
rect 1074 414 1134 463
rect 1074 380 1087 414
rect 1121 380 1134 414
rect 1074 368 1134 380
rect 1164 572 1224 592
rect 1164 538 1177 572
rect 1211 538 1224 572
rect 1164 478 1224 538
rect 1164 444 1177 478
rect 1211 444 1224 478
rect 1164 368 1224 444
rect 1254 580 1314 592
rect 1254 546 1267 580
rect 1301 546 1314 580
rect 1254 497 1314 546
rect 1254 463 1267 497
rect 1301 463 1314 497
rect 1254 414 1314 463
rect 1254 380 1267 414
rect 1301 380 1314 414
rect 1254 368 1314 380
rect 1344 580 1400 592
rect 1344 546 1358 580
rect 1392 546 1400 580
rect 1344 510 1400 546
rect 1344 476 1358 510
rect 1392 476 1400 510
rect 1344 440 1400 476
rect 1344 406 1358 440
rect 1392 406 1400 440
rect 1344 368 1400 406
<< ndiffc >>
rect 39 150 73 184
rect 141 118 175 152
rect 241 176 275 210
rect 241 86 275 120
rect 353 176 387 210
rect 353 86 387 120
rect 439 92 473 126
rect 525 176 559 210
rect 611 92 645 126
rect 711 176 745 210
rect 711 86 745 120
rect 811 92 845 126
rect 897 176 931 210
rect 983 92 1017 126
rect 1075 176 1109 210
rect 1167 92 1201 126
rect 1267 176 1301 210
rect 1267 86 1301 120
rect 1367 170 1401 204
rect 1367 86 1401 120
<< pdiffc >>
rect 39 490 73 524
rect 39 395 73 429
rect 131 490 165 524
rect 234 546 268 580
rect 234 463 268 497
rect 234 380 268 414
rect 346 546 380 580
rect 346 463 380 497
rect 346 380 380 414
rect 436 546 470 580
rect 436 448 470 482
rect 526 546 560 580
rect 526 463 560 497
rect 526 380 560 414
rect 626 546 660 580
rect 626 463 660 497
rect 626 380 660 414
rect 726 546 760 580
rect 726 463 760 497
rect 726 380 760 414
rect 816 546 850 580
rect 816 444 850 478
rect 906 546 940 580
rect 906 463 940 497
rect 906 380 940 414
rect 996 546 1030 580
rect 996 444 1030 478
rect 1087 546 1121 580
rect 1087 463 1121 497
rect 1087 380 1121 414
rect 1177 538 1211 572
rect 1177 444 1211 478
rect 1267 546 1301 580
rect 1267 463 1301 497
rect 1267 380 1301 414
rect 1358 546 1392 580
rect 1358 476 1392 510
rect 1358 406 1392 440
<< poly >>
rect 191 592 221 618
rect 393 592 423 618
rect 483 592 513 618
rect 573 592 603 618
rect 673 592 703 618
rect 773 592 803 618
rect 863 592 893 618
rect 953 592 983 618
rect 1044 592 1074 618
rect 1134 592 1164 618
rect 1224 592 1254 618
rect 1314 592 1344 618
rect 86 536 116 562
rect 86 353 116 368
rect 191 353 221 368
rect 393 353 423 368
rect 483 353 513 368
rect 573 353 603 368
rect 673 353 703 368
rect 773 353 803 368
rect 863 353 893 368
rect 953 353 983 368
rect 1044 353 1074 368
rect 1134 353 1164 368
rect 1224 353 1254 368
rect 1314 353 1344 368
rect 83 336 116 353
rect 48 320 114 336
rect 188 326 224 353
rect 390 326 426 353
rect 480 326 516 353
rect 570 326 606 353
rect 48 286 64 320
rect 98 286 114 320
rect 48 270 114 286
rect 84 222 114 270
rect 162 310 230 326
rect 162 276 178 310
rect 212 276 230 310
rect 162 260 230 276
rect 305 310 606 326
rect 305 276 321 310
rect 355 276 389 310
rect 423 276 457 310
rect 491 276 606 310
rect 305 260 606 276
rect 670 326 706 353
rect 770 326 806 353
rect 860 326 896 353
rect 950 326 986 353
rect 1041 326 1077 353
rect 1131 326 1167 353
rect 1221 326 1257 353
rect 1311 326 1347 353
rect 670 310 1347 326
rect 670 276 686 310
rect 720 276 754 310
rect 788 276 822 310
rect 856 276 890 310
rect 924 276 958 310
rect 992 276 1026 310
rect 1060 276 1094 310
rect 1128 276 1162 310
rect 1196 276 1347 310
rect 670 260 1347 276
rect 200 222 230 260
rect 398 222 428 260
rect 484 222 514 260
rect 570 222 600 260
rect 670 222 700 260
rect 756 222 786 260
rect 856 222 886 260
rect 942 222 972 260
rect 1028 222 1058 260
rect 1126 222 1156 260
rect 1226 222 1256 260
rect 1312 222 1342 260
rect 84 86 114 112
rect 200 48 230 74
rect 398 48 428 74
rect 484 48 514 74
rect 570 48 600 74
rect 670 48 700 74
rect 756 48 786 74
rect 856 48 886 74
rect 942 48 972 74
rect 1028 48 1058 74
rect 1126 48 1156 74
rect 1226 48 1256 74
rect 1312 48 1342 74
<< polycont >>
rect 64 286 98 320
rect 178 276 212 310
rect 321 276 355 310
rect 389 276 423 310
rect 457 276 491 310
rect 686 276 720 310
rect 754 276 788 310
rect 822 276 856 310
rect 890 276 924 310
rect 958 276 992 310
rect 1026 276 1060 310
rect 1094 276 1128 310
rect 1162 276 1196 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 524 76 540
rect 23 490 39 524
rect 73 490 76 524
rect 23 440 76 490
rect 113 524 184 649
rect 113 490 131 524
rect 165 490 184 524
rect 113 474 184 490
rect 218 580 296 596
rect 218 546 234 580
rect 268 546 296 580
rect 218 497 296 546
rect 218 463 234 497
rect 268 463 296 497
rect 23 429 184 440
rect 23 395 39 429
rect 73 395 184 429
rect 23 390 184 395
rect 25 320 114 356
rect 25 286 64 320
rect 98 286 114 320
rect 25 270 114 286
rect 150 326 184 390
rect 218 414 296 463
rect 218 380 234 414
rect 268 380 296 414
rect 218 364 296 380
rect 330 580 396 596
rect 330 546 346 580
rect 380 546 396 580
rect 330 497 396 546
rect 330 463 346 497
rect 380 463 396 497
rect 330 414 396 463
rect 430 580 476 649
rect 430 546 436 580
rect 470 546 476 580
rect 430 482 476 546
rect 430 448 436 482
rect 470 448 476 482
rect 430 432 476 448
rect 510 580 576 596
rect 510 546 526 580
rect 560 546 576 580
rect 510 497 576 546
rect 510 463 526 497
rect 560 463 576 497
rect 330 380 346 414
rect 380 398 396 414
rect 510 414 576 463
rect 510 398 526 414
rect 380 380 526 398
rect 560 380 576 414
rect 330 364 576 380
rect 610 580 676 649
rect 610 546 626 580
rect 660 546 676 580
rect 610 497 676 546
rect 610 463 626 497
rect 660 463 676 497
rect 610 414 676 463
rect 610 380 626 414
rect 660 380 676 414
rect 610 364 676 380
rect 713 580 766 596
rect 713 546 726 580
rect 760 546 766 580
rect 713 497 766 546
rect 713 463 726 497
rect 760 463 766 497
rect 713 414 766 463
rect 807 580 858 649
rect 807 546 816 580
rect 850 546 858 580
rect 807 478 858 546
rect 807 444 816 478
rect 850 444 858 478
rect 807 428 858 444
rect 899 580 949 596
rect 899 546 906 580
rect 940 546 949 580
rect 899 497 949 546
rect 899 463 906 497
rect 940 463 949 497
rect 713 380 726 414
rect 760 394 766 414
rect 899 414 949 463
rect 986 580 1041 649
rect 986 546 996 580
rect 1030 546 1041 580
rect 986 478 1041 546
rect 986 444 996 478
rect 1030 444 1041 478
rect 986 428 1041 444
rect 1077 580 1131 596
rect 1077 546 1087 580
rect 1121 546 1131 580
rect 1077 497 1131 546
rect 1077 463 1087 497
rect 1121 463 1131 497
rect 899 394 906 414
rect 760 380 906 394
rect 940 394 949 414
rect 1077 414 1131 463
rect 1167 572 1221 649
rect 1167 538 1177 572
rect 1211 538 1221 572
rect 1167 478 1221 538
rect 1167 444 1177 478
rect 1211 444 1221 478
rect 1167 428 1221 444
rect 1257 580 1311 596
rect 1257 546 1267 580
rect 1301 546 1311 580
rect 1257 497 1311 546
rect 1257 463 1267 497
rect 1301 463 1311 497
rect 1077 394 1087 414
rect 940 380 1087 394
rect 1121 394 1131 414
rect 1257 414 1311 463
rect 1257 394 1267 414
rect 1121 380 1267 394
rect 1301 380 1311 414
rect 1347 580 1408 649
rect 1347 546 1358 580
rect 1392 546 1408 580
rect 1347 510 1408 546
rect 1347 476 1358 510
rect 1392 476 1408 510
rect 1347 440 1408 476
rect 1347 406 1358 440
rect 1392 406 1408 440
rect 1347 390 1408 406
rect 262 326 296 364
rect 534 326 576 364
rect 713 360 1311 380
rect 1251 356 1311 360
rect 150 310 228 326
rect 150 276 178 310
rect 212 276 228 310
rect 150 260 228 276
rect 262 310 500 326
rect 262 276 321 310
rect 355 276 389 310
rect 423 276 457 310
rect 491 276 500 310
rect 262 260 500 276
rect 534 310 1204 326
rect 534 276 686 310
rect 720 276 754 310
rect 788 276 822 310
rect 856 276 890 310
rect 924 276 958 310
rect 992 276 1026 310
rect 1060 276 1094 310
rect 1128 276 1162 310
rect 1196 276 1204 310
rect 534 260 1204 276
rect 150 236 184 260
rect 23 202 184 236
rect 262 226 296 260
rect 534 226 625 260
rect 1251 254 1415 356
rect 1251 226 1317 254
rect 225 210 296 226
rect 23 184 89 202
rect 23 150 39 184
rect 73 150 89 184
rect 225 176 241 210
rect 275 176 296 210
rect 23 108 89 150
rect 125 152 191 168
rect 125 118 141 152
rect 175 118 191 152
rect 125 17 191 118
rect 225 120 296 176
rect 225 86 241 120
rect 275 86 296 120
rect 225 70 296 86
rect 337 210 625 226
rect 337 176 353 210
rect 387 176 525 210
rect 559 176 625 210
rect 695 210 1317 226
rect 695 176 711 210
rect 745 176 897 210
rect 931 176 1075 210
rect 1109 176 1267 210
rect 1301 176 1317 210
rect 337 120 387 176
rect 337 86 353 120
rect 337 70 387 86
rect 423 126 489 142
rect 423 92 439 126
rect 473 92 489 126
rect 423 17 489 92
rect 595 126 661 142
rect 595 92 611 126
rect 645 92 661 126
rect 595 17 661 92
rect 695 120 761 176
rect 695 86 711 120
rect 745 86 761 120
rect 695 70 761 86
rect 795 126 861 142
rect 795 92 811 126
rect 845 92 861 126
rect 795 17 861 92
rect 967 126 1033 142
rect 967 92 983 126
rect 1017 92 1033 126
rect 967 17 1033 92
rect 1151 126 1217 142
rect 1151 92 1167 126
rect 1201 92 1217 126
rect 1151 17 1217 92
rect 1251 120 1317 176
rect 1251 86 1267 120
rect 1301 86 1317 120
rect 1251 70 1317 86
rect 1351 204 1417 220
rect 1351 170 1367 204
rect 1401 170 1417 204
rect 1351 120 1417 170
rect 1351 86 1367 120
rect 1401 86 1417 120
rect 1351 17 1417 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 bufbuf_8
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3943392
string GDS_START 3932438
<< end >>
