magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
rect 749 325 2412 331
rect 749 311 2066 325
<< pwell >>
rect 1134 235 1485 265
rect 1884 235 2159 265
rect 46 176 705 235
rect 1134 179 2159 235
rect 1134 176 2783 179
rect 46 49 2783 176
rect 0 0 2784 49
<< scnmos >>
rect 129 125 159 209
rect 207 125 237 209
rect 321 125 351 209
rect 399 125 429 209
rect 501 125 531 209
rect 593 125 623 209
rect 1233 155 1263 239
rect 1373 155 1403 239
rect 790 66 820 150
rect 862 66 892 150
rect 948 66 978 150
rect 1020 66 1050 150
rect 1576 125 1606 209
rect 1692 125 1722 209
rect 1764 125 1794 209
rect 1963 155 1993 239
rect 2049 155 2079 239
rect 2243 69 2273 153
rect 2329 69 2359 153
rect 2401 69 2431 153
rect 2598 69 2628 153
rect 2670 69 2700 153
<< scpmoshvt >>
rect 84 409 134 609
rect 301 417 351 617
rect 407 417 457 617
rect 501 417 551 617
rect 607 417 657 617
rect 842 347 892 547
rect 948 347 998 547
rect 1372 347 1422 547
rect 1478 347 1528 547
rect 1576 347 1626 547
rect 1767 347 1817 547
rect 1907 347 1957 547
rect 2045 361 2095 561
rect 2148 361 2198 561
rect 2269 361 2319 561
rect 2650 388 2700 588
<< ndiff >>
rect 72 184 129 209
rect 72 150 84 184
rect 118 150 129 184
rect 72 125 129 150
rect 159 125 207 209
rect 237 176 321 209
rect 237 142 248 176
rect 282 142 321 176
rect 237 125 321 142
rect 351 125 399 209
rect 429 181 501 209
rect 429 147 456 181
rect 490 147 501 181
rect 429 125 501 147
rect 531 125 593 209
rect 623 184 679 209
rect 623 150 634 184
rect 668 150 679 184
rect 1160 205 1233 239
rect 1160 171 1172 205
rect 1206 171 1233 205
rect 1160 155 1233 171
rect 1263 227 1373 239
rect 1263 193 1328 227
rect 1362 193 1373 227
rect 1263 155 1373 193
rect 1403 211 1459 239
rect 1403 177 1414 211
rect 1448 177 1459 211
rect 1403 155 1459 177
rect 623 125 679 150
rect 733 125 790 150
rect 733 91 745 125
rect 779 91 790 125
rect 733 66 790 91
rect 820 66 862 150
rect 892 113 948 150
rect 892 79 903 113
rect 937 79 948 113
rect 892 66 948 79
rect 978 66 1020 150
rect 1050 125 1106 150
rect 1050 91 1061 125
rect 1095 91 1106 125
rect 1050 66 1106 91
rect 1519 175 1576 209
rect 1519 141 1531 175
rect 1565 141 1576 175
rect 1519 125 1576 141
rect 1606 127 1692 209
rect 1606 125 1632 127
rect 1621 93 1632 125
rect 1666 125 1692 127
rect 1722 125 1764 209
rect 1794 184 1850 209
rect 1794 150 1805 184
rect 1839 150 1850 184
rect 1794 125 1850 150
rect 1666 93 1677 125
rect 1621 81 1677 93
rect 1910 214 1963 239
rect 1910 180 1918 214
rect 1952 180 1963 214
rect 1910 155 1963 180
rect 1993 227 2049 239
rect 1993 193 2004 227
rect 2038 193 2049 227
rect 1993 155 2049 193
rect 2079 155 2133 239
rect 2094 99 2133 155
rect 2075 87 2133 99
rect 2075 53 2087 87
rect 2121 53 2133 87
rect 2187 128 2243 153
rect 2187 94 2198 128
rect 2232 94 2243 128
rect 2187 69 2243 94
rect 2273 128 2329 153
rect 2273 94 2284 128
rect 2318 94 2329 128
rect 2273 69 2329 94
rect 2359 69 2401 153
rect 2431 128 2487 153
rect 2431 94 2442 128
rect 2476 94 2487 128
rect 2431 69 2487 94
rect 2541 128 2598 153
rect 2541 94 2553 128
rect 2587 94 2598 128
rect 2541 69 2598 94
rect 2628 69 2670 153
rect 2700 128 2757 153
rect 2700 94 2711 128
rect 2745 94 2757 128
rect 2700 69 2757 94
rect 2075 41 2133 53
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 190 609
rect 134 563 145 597
rect 179 563 190 597
rect 134 526 190 563
rect 134 492 145 526
rect 179 492 190 526
rect 134 455 190 492
rect 134 421 145 455
rect 179 421 190 455
rect 134 409 190 421
rect 244 597 301 617
rect 244 563 256 597
rect 290 563 301 597
rect 244 463 301 563
rect 244 429 256 463
rect 290 429 301 463
rect 244 417 301 429
rect 351 464 407 617
rect 351 430 362 464
rect 396 430 407 464
rect 351 417 407 430
rect 457 417 501 617
rect 551 605 607 617
rect 551 571 562 605
rect 596 571 607 605
rect 551 417 607 571
rect 657 574 714 617
rect 657 540 668 574
rect 702 540 714 574
rect 657 417 714 540
rect 785 394 842 547
rect 785 360 797 394
rect 831 360 842 394
rect 785 347 842 360
rect 892 535 948 547
rect 892 501 903 535
rect 937 501 948 535
rect 892 347 948 501
rect 998 394 1055 547
rect 2593 576 2650 588
rect 1972 549 2045 561
rect 1972 547 1984 549
rect 998 360 1009 394
rect 1043 360 1055 394
rect 998 347 1055 360
rect 1315 535 1372 547
rect 1315 501 1327 535
rect 1361 501 1372 535
rect 1315 464 1372 501
rect 1315 430 1327 464
rect 1361 430 1372 464
rect 1315 393 1372 430
rect 1315 359 1327 393
rect 1361 359 1372 393
rect 1315 347 1372 359
rect 1422 535 1478 547
rect 1422 501 1433 535
rect 1467 501 1478 535
rect 1422 464 1478 501
rect 1422 430 1433 464
rect 1467 430 1478 464
rect 1422 393 1478 430
rect 1422 359 1433 393
rect 1467 359 1478 393
rect 1422 347 1478 359
rect 1528 347 1576 547
rect 1626 535 1767 547
rect 1626 501 1637 535
rect 1671 501 1767 535
rect 1626 453 1767 501
rect 1626 419 1637 453
rect 1671 419 1767 453
rect 1626 347 1767 419
rect 1817 535 1907 547
rect 1817 501 1837 535
rect 1871 501 1907 535
rect 1817 464 1907 501
rect 1817 430 1837 464
rect 1871 430 1907 464
rect 1817 393 1907 430
rect 1817 359 1837 393
rect 1871 359 1907 393
rect 1817 347 1907 359
rect 1957 515 1984 547
rect 2018 515 2045 549
rect 1957 471 2045 515
rect 1957 437 1984 471
rect 2018 437 2045 471
rect 1957 393 2045 437
rect 1957 359 1984 393
rect 2018 361 2045 393
rect 2095 361 2148 561
rect 2198 549 2269 561
rect 2198 515 2209 549
rect 2243 515 2269 549
rect 2198 415 2269 515
rect 2198 381 2209 415
rect 2243 381 2269 415
rect 2198 361 2269 381
rect 2319 549 2376 561
rect 2319 515 2330 549
rect 2364 515 2376 549
rect 2319 415 2376 515
rect 2319 381 2330 415
rect 2364 381 2376 415
rect 2593 542 2605 576
rect 2639 542 2650 576
rect 2593 505 2650 542
rect 2593 471 2605 505
rect 2639 471 2650 505
rect 2593 434 2650 471
rect 2593 400 2605 434
rect 2639 400 2650 434
rect 2593 388 2650 400
rect 2700 576 2757 588
rect 2700 542 2711 576
rect 2745 542 2757 576
rect 2700 505 2757 542
rect 2700 471 2711 505
rect 2745 471 2757 505
rect 2700 434 2757 471
rect 2700 400 2711 434
rect 2745 400 2757 434
rect 2700 388 2757 400
rect 2319 361 2376 381
rect 2018 359 2030 361
rect 1957 347 2030 359
<< ndiffc >>
rect 84 150 118 184
rect 248 142 282 176
rect 456 147 490 181
rect 634 150 668 184
rect 1172 171 1206 205
rect 1328 193 1362 227
rect 1414 177 1448 211
rect 745 91 779 125
rect 903 79 937 113
rect 1061 91 1095 125
rect 1531 141 1565 175
rect 1632 93 1666 127
rect 1805 150 1839 184
rect 1918 180 1952 214
rect 2004 193 2038 227
rect 2087 53 2121 87
rect 2198 94 2232 128
rect 2284 94 2318 128
rect 2442 94 2476 128
rect 2553 94 2587 128
rect 2711 94 2745 128
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 256 563 290 597
rect 256 429 290 463
rect 362 430 396 464
rect 562 571 596 605
rect 668 540 702 574
rect 797 360 831 394
rect 903 501 937 535
rect 1009 360 1043 394
rect 1327 501 1361 535
rect 1327 430 1361 464
rect 1327 359 1361 393
rect 1433 501 1467 535
rect 1433 430 1467 464
rect 1433 359 1467 393
rect 1637 501 1671 535
rect 1637 419 1671 453
rect 1837 501 1871 535
rect 1837 430 1871 464
rect 1837 359 1871 393
rect 1984 515 2018 549
rect 1984 437 2018 471
rect 1984 359 2018 393
rect 2209 515 2243 549
rect 2209 381 2243 415
rect 2330 515 2364 549
rect 2330 381 2364 415
rect 2605 542 2639 576
rect 2605 471 2639 505
rect 2605 400 2639 434
rect 2711 542 2745 576
rect 2711 471 2745 505
rect 2711 400 2745 434
<< poly >>
rect 84 609 134 635
rect 301 617 351 643
rect 407 617 457 643
rect 501 617 551 643
rect 607 617 657 643
rect 1134 615 2095 645
rect 842 547 892 573
rect 948 547 998 573
rect 84 369 134 409
rect 84 353 175 369
rect 301 367 351 417
rect 407 377 457 417
rect 84 319 125 353
rect 159 333 175 353
rect 285 351 351 367
rect 159 319 237 333
rect 84 303 237 319
rect 129 209 159 303
rect 207 209 237 303
rect 285 317 301 351
rect 335 317 351 351
rect 285 283 351 317
rect 285 249 301 283
rect 335 249 351 283
rect 285 233 351 249
rect 393 361 459 377
rect 393 327 409 361
rect 443 327 459 361
rect 393 293 459 327
rect 393 259 409 293
rect 443 259 459 293
rect 393 243 459 259
rect 321 209 351 233
rect 399 209 429 243
rect 501 224 551 417
rect 607 383 657 417
rect 593 367 667 383
rect 593 333 617 367
rect 651 333 667 367
rect 1134 395 1164 615
rect 1372 547 1422 615
rect 1478 547 1528 573
rect 1576 547 1626 573
rect 1767 547 1817 573
rect 1907 547 1957 573
rect 2045 561 2095 615
rect 2650 588 2700 614
rect 2148 561 2198 587
rect 2269 561 2319 587
rect 1098 379 1164 395
rect 593 299 667 333
rect 842 302 892 347
rect 948 306 998 347
rect 1098 345 1114 379
rect 1148 345 1164 379
rect 1098 311 1164 345
rect 1372 321 1422 347
rect 593 265 617 299
rect 651 265 667 299
rect 593 249 667 265
rect 790 286 892 302
rect 790 252 806 286
rect 840 252 892 286
rect 501 209 531 224
rect 593 209 623 249
rect 790 236 892 252
rect 790 150 820 236
rect 862 150 892 236
rect 943 290 1009 306
rect 943 256 959 290
rect 993 256 1009 290
rect 1098 277 1114 311
rect 1148 291 1164 311
rect 1148 277 1263 291
rect 1098 261 1263 277
rect 943 222 1009 256
rect 1233 239 1263 261
rect 1373 239 1403 265
rect 1478 254 1528 347
rect 943 188 959 222
rect 993 202 1009 222
rect 993 188 1050 202
rect 943 172 1050 188
rect 948 150 978 172
rect 1020 150 1050 172
rect 1474 224 1528 254
rect 1576 297 1626 347
rect 1767 315 1817 347
rect 1692 299 1817 315
rect 1576 281 1642 297
rect 1576 247 1592 281
rect 1626 247 1642 281
rect 1576 231 1642 247
rect 1692 265 1708 299
rect 1742 265 1817 299
rect 1907 284 1957 347
rect 2045 335 2095 361
rect 2049 330 2095 335
rect 1692 249 1817 265
rect 1865 254 1993 284
rect 129 99 159 125
rect 207 51 237 125
rect 321 99 351 125
rect 399 99 429 125
rect 501 51 531 125
rect 593 99 623 125
rect 1233 129 1263 155
rect 207 21 531 51
rect 790 40 820 66
rect 862 40 892 66
rect 948 40 978 66
rect 1020 51 1050 66
rect 1373 51 1403 155
rect 1474 51 1504 224
rect 1576 209 1606 231
rect 1692 209 1722 249
rect 1764 209 1794 249
rect 1576 99 1606 125
rect 1692 99 1722 125
rect 1764 99 1794 125
rect 1865 51 1895 254
rect 1963 239 1993 254
rect 2049 239 2079 330
rect 2148 259 2198 361
rect 2269 329 2319 361
rect 2269 313 2359 329
rect 2269 279 2285 313
rect 2319 279 2359 313
rect 2269 263 2359 279
rect 2479 311 2545 327
rect 2479 277 2495 311
rect 2529 277 2545 311
rect 2148 243 2221 259
rect 2148 209 2171 243
rect 2205 215 2221 243
rect 2329 233 2431 263
rect 2205 209 2273 215
rect 2148 185 2273 209
rect 1963 129 1993 155
rect 2049 129 2079 155
rect 2243 153 2273 185
rect 2329 153 2359 233
rect 2401 153 2431 233
rect 2479 243 2545 277
rect 2479 209 2495 243
rect 2529 223 2545 243
rect 2650 223 2700 388
rect 2529 209 2700 223
rect 2479 193 2700 209
rect 2598 153 2628 193
rect 2670 153 2700 193
rect 1020 21 1895 51
rect 2243 43 2273 69
rect 2329 43 2359 69
rect 2401 43 2431 69
rect 2598 43 2628 69
rect 2670 43 2700 69
<< polycont >>
rect 125 319 159 353
rect 301 317 335 351
rect 301 249 335 283
rect 409 327 443 361
rect 409 259 443 293
rect 617 333 651 367
rect 1114 345 1148 379
rect 617 265 651 299
rect 806 252 840 286
rect 959 256 993 290
rect 1114 277 1148 311
rect 959 188 993 222
rect 1592 247 1626 281
rect 1708 265 1742 299
rect 2285 279 2319 313
rect 2495 277 2529 311
rect 2171 209 2205 243
rect 2495 209 2529 243
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 597 73 613
rect 23 563 39 597
rect 23 526 73 563
rect 23 492 39 526
rect 23 455 73 492
rect 23 421 39 455
rect 23 267 73 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 240 597 306 613
rect 240 563 256 597
rect 290 563 306 597
rect 546 605 612 649
rect 546 571 562 605
rect 596 571 612 605
rect 652 574 718 613
rect 240 535 306 563
rect 652 540 668 574
rect 702 540 718 574
rect 652 535 718 540
rect 240 501 718 535
rect 887 535 953 649
rect 887 501 903 535
rect 937 501 953 535
rect 1311 535 1377 551
rect 1311 501 1327 535
rect 1361 501 1377 535
rect 240 463 306 501
rect 1311 465 1377 501
rect 240 429 256 463
rect 290 429 306 463
rect 240 413 306 429
rect 346 464 1377 465
rect 346 430 362 464
rect 396 431 1327 464
rect 396 430 529 431
rect 346 413 529 430
rect 109 353 175 369
rect 109 319 125 353
rect 159 319 175 353
rect 109 303 175 319
rect 285 351 351 367
rect 285 317 301 351
rect 335 317 351 351
rect 285 283 351 317
rect 285 267 301 283
rect 23 249 301 267
rect 335 249 351 283
rect 23 233 351 249
rect 393 361 459 377
rect 393 327 409 361
rect 443 327 459 361
rect 393 293 459 327
rect 393 259 409 293
rect 443 259 459 293
rect 393 243 459 259
rect 23 184 134 233
rect 495 207 529 413
rect 1242 430 1327 431
rect 1361 430 1377 464
rect 781 394 926 395
rect 601 367 743 383
rect 601 333 617 367
rect 651 333 743 367
rect 781 360 797 394
rect 831 360 926 394
rect 781 343 926 360
rect 993 394 1164 395
rect 993 360 1009 394
rect 1043 379 1164 394
rect 1043 360 1114 379
rect 993 345 1114 360
rect 1148 345 1164 379
rect 993 343 1164 345
rect 601 299 743 333
rect 892 306 926 343
rect 1045 311 1164 343
rect 601 265 617 299
rect 651 265 743 299
rect 601 249 743 265
rect 790 286 856 302
rect 790 252 806 286
rect 840 252 856 286
rect 790 236 856 252
rect 892 290 1009 306
rect 892 256 959 290
rect 993 256 1009 290
rect 892 222 1009 256
rect 23 150 84 184
rect 118 150 134 184
rect 23 121 134 150
rect 232 176 298 197
rect 232 142 248 176
rect 282 142 298 176
rect 232 17 298 142
rect 440 181 529 207
rect 440 147 456 181
rect 490 147 529 181
rect 440 121 529 147
rect 618 184 684 213
rect 892 200 959 222
rect 618 150 634 184
rect 668 150 684 184
rect 618 17 684 150
rect 729 188 959 200
rect 993 188 1009 222
rect 729 166 1009 188
rect 1045 277 1114 311
rect 1148 277 1164 311
rect 1045 261 1164 277
rect 1242 393 1377 430
rect 1242 359 1327 393
rect 1361 359 1377 393
rect 1242 343 1377 359
rect 1417 535 1483 551
rect 1417 501 1433 535
rect 1467 501 1483 535
rect 1417 464 1483 501
rect 1417 430 1433 464
rect 1467 430 1483 464
rect 1417 393 1483 430
rect 1621 535 1687 649
rect 1621 501 1637 535
rect 1671 501 1687 535
rect 1621 453 1687 501
rect 1621 419 1637 453
rect 1671 419 1687 453
rect 1621 403 1687 419
rect 1821 535 1887 551
rect 1821 501 1837 535
rect 1871 501 1887 535
rect 1821 464 1887 501
rect 1821 430 1837 464
rect 1871 430 1887 464
rect 1417 359 1433 393
rect 1467 367 1483 393
rect 1821 393 1887 430
rect 1467 359 1758 367
rect 729 125 795 166
rect 729 91 745 125
rect 779 91 795 125
rect 729 62 795 91
rect 887 113 953 130
rect 887 79 903 113
rect 937 79 953 113
rect 887 17 953 79
rect 1045 125 1111 261
rect 1045 91 1061 125
rect 1095 91 1111 125
rect 1045 62 1111 91
rect 1156 205 1206 225
rect 1156 171 1172 205
rect 1156 87 1206 171
rect 1242 157 1276 343
rect 1417 333 1758 359
rect 1417 307 1483 333
rect 1312 273 1483 307
rect 1692 299 1758 333
rect 1576 281 1642 297
rect 1312 227 1378 273
rect 1576 247 1592 281
rect 1626 247 1642 281
rect 1692 265 1708 299
rect 1742 265 1758 299
rect 1692 249 1758 265
rect 1821 359 1837 393
rect 1871 359 1887 393
rect 1821 343 1887 359
rect 1968 549 2034 565
rect 1968 515 1984 549
rect 2018 515 2034 549
rect 1968 471 2034 515
rect 1968 437 1984 471
rect 2018 437 2034 471
rect 1968 393 2034 437
rect 1968 359 1984 393
rect 2018 359 2034 393
rect 2193 549 2259 649
rect 2521 576 2655 592
rect 2193 515 2209 549
rect 2243 515 2259 549
rect 2193 415 2259 515
rect 2193 381 2209 415
rect 2243 381 2259 415
rect 2193 365 2259 381
rect 2314 549 2405 565
rect 2314 515 2330 549
rect 2364 515 2405 549
rect 2314 415 2405 515
rect 2314 381 2330 415
rect 2364 381 2405 415
rect 2521 542 2605 576
rect 2639 542 2655 576
rect 2521 505 2655 542
rect 2521 471 2605 505
rect 2639 471 2655 505
rect 2521 434 2655 471
rect 2521 400 2605 434
rect 2639 400 2655 434
rect 2521 384 2655 400
rect 2695 576 2761 649
rect 2695 542 2711 576
rect 2745 542 2761 576
rect 2695 505 2761 542
rect 2695 471 2711 505
rect 2745 471 2761 505
rect 2695 434 2761 471
rect 2695 400 2711 434
rect 2745 400 2761 434
rect 2695 384 2761 400
rect 2314 365 2405 381
rect 1312 193 1328 227
rect 1362 193 1378 227
rect 1414 211 1464 237
rect 1576 231 1642 247
rect 1448 177 1464 211
rect 1608 213 1642 231
rect 1821 213 1855 343
rect 1968 329 2034 359
rect 1968 313 2335 329
rect 1968 295 2285 313
rect 1414 157 1464 177
rect 1242 123 1464 157
rect 1515 175 1565 195
rect 1608 184 1855 213
rect 1608 179 1805 184
rect 1515 141 1531 175
rect 1789 150 1805 179
rect 1839 150 1855 184
rect 1515 87 1565 141
rect 1156 53 1565 87
rect 1616 127 1682 143
rect 1616 93 1632 127
rect 1666 93 1682 127
rect 1616 17 1682 93
rect 1789 87 1855 150
rect 1906 214 1954 243
rect 1906 180 1918 214
rect 1952 180 1954 214
rect 1988 227 2054 295
rect 2269 279 2285 295
rect 2319 279 2335 313
rect 2269 263 2335 279
rect 1988 193 2004 227
rect 2038 193 2054 227
rect 2155 243 2221 259
rect 2155 209 2171 243
rect 2205 227 2221 243
rect 2371 227 2405 365
rect 2479 311 2545 327
rect 2479 277 2495 311
rect 2529 277 2545 311
rect 2479 243 2545 277
rect 2479 227 2495 243
rect 2205 209 2495 227
rect 2529 209 2545 243
rect 2155 193 2545 209
rect 1906 157 1954 180
rect 2426 157 2460 193
rect 2581 157 2615 384
rect 1906 128 2232 157
rect 1906 123 2198 128
rect 2182 94 2198 123
rect 1789 53 2087 87
rect 2121 53 2137 87
rect 2182 65 2232 94
rect 2268 128 2334 157
rect 2268 94 2284 128
rect 2318 94 2334 128
rect 2268 17 2334 94
rect 2426 128 2492 157
rect 2426 94 2442 128
rect 2476 94 2492 128
rect 2426 65 2492 94
rect 2537 128 2615 157
rect 2537 94 2553 128
rect 2587 94 2615 128
rect 2537 65 2615 94
rect 2695 128 2761 157
rect 2695 94 2711 128
rect 2745 94 2761 128
rect 2695 17 2761 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxtp_lp
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2527 464 2561 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2527 538 2561 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4019450
string GDS_START 4002594
<< end >>
