magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 93 49 2015 241
rect 0 0 2016 49
<< scnmos >>
rect 172 47 202 215
rect 258 47 288 215
rect 344 47 374 215
rect 430 47 460 215
rect 516 47 546 215
rect 602 47 632 215
rect 688 47 718 215
rect 830 47 860 215
rect 916 47 946 215
rect 1002 47 1032 215
rect 1088 47 1118 215
rect 1202 47 1232 215
rect 1304 47 1334 215
rect 1390 47 1420 215
rect 1476 47 1506 215
rect 1562 47 1592 215
rect 1648 47 1678 215
rect 1734 47 1764 215
rect 1820 47 1850 215
rect 1906 47 1936 215
<< scpmoshvt >>
rect 138 367 168 619
rect 224 367 254 619
rect 310 367 340 619
rect 396 367 426 619
rect 586 367 616 619
rect 672 367 702 619
rect 758 367 788 619
rect 844 367 874 619
rect 930 367 960 619
rect 1016 367 1046 619
rect 1102 367 1132 619
rect 1188 367 1218 619
rect 1298 367 1328 619
rect 1390 367 1420 619
rect 1476 367 1506 619
rect 1562 367 1592 619
rect 1648 367 1678 619
rect 1734 367 1764 619
rect 1820 367 1850 619
rect 1906 367 1936 619
<< ndiff >>
rect 119 203 172 215
rect 119 169 127 203
rect 161 169 172 203
rect 119 93 172 169
rect 119 59 127 93
rect 161 59 172 93
rect 119 47 172 59
rect 202 192 258 215
rect 202 158 213 192
rect 247 158 258 192
rect 202 101 258 158
rect 202 67 213 101
rect 247 67 258 101
rect 202 47 258 67
rect 288 132 344 215
rect 288 98 299 132
rect 333 98 344 132
rect 288 47 344 98
rect 374 192 430 215
rect 374 158 385 192
rect 419 158 430 192
rect 374 101 430 158
rect 374 67 385 101
rect 419 67 430 101
rect 374 47 430 67
rect 460 132 516 215
rect 460 98 471 132
rect 505 98 516 132
rect 460 47 516 98
rect 546 151 602 215
rect 546 117 557 151
rect 591 117 602 151
rect 546 47 602 117
rect 632 93 688 215
rect 632 59 643 93
rect 677 59 688 93
rect 632 47 688 59
rect 718 101 830 215
rect 718 67 729 101
rect 763 67 830 101
rect 718 47 830 67
rect 860 202 916 215
rect 860 168 871 202
rect 905 168 916 202
rect 860 47 916 168
rect 946 101 1002 215
rect 946 67 957 101
rect 991 67 1002 101
rect 946 47 1002 67
rect 1032 202 1088 215
rect 1032 168 1043 202
rect 1077 168 1088 202
rect 1032 47 1088 168
rect 1118 101 1202 215
rect 1118 67 1157 101
rect 1191 67 1202 101
rect 1118 47 1202 67
rect 1232 130 1304 215
rect 1232 96 1243 130
rect 1277 96 1304 130
rect 1232 47 1304 96
rect 1334 93 1390 215
rect 1334 59 1345 93
rect 1379 59 1390 93
rect 1334 47 1390 59
rect 1420 190 1476 215
rect 1420 156 1431 190
rect 1465 156 1476 190
rect 1420 47 1476 156
rect 1506 93 1562 215
rect 1506 59 1517 93
rect 1551 59 1562 93
rect 1506 47 1562 59
rect 1592 190 1648 215
rect 1592 156 1603 190
rect 1637 156 1648 190
rect 1592 47 1648 156
rect 1678 192 1734 215
rect 1678 158 1689 192
rect 1723 158 1734 192
rect 1678 101 1734 158
rect 1678 67 1689 101
rect 1723 67 1734 101
rect 1678 47 1734 67
rect 1764 132 1820 215
rect 1764 98 1775 132
rect 1809 98 1820 132
rect 1764 47 1820 98
rect 1850 192 1906 215
rect 1850 158 1861 192
rect 1895 158 1906 192
rect 1850 101 1906 158
rect 1850 67 1861 101
rect 1895 67 1906 101
rect 1850 47 1906 67
rect 1936 203 1989 215
rect 1936 169 1947 203
rect 1981 169 1989 203
rect 1936 93 1989 169
rect 1936 59 1947 93
rect 1981 59 1989 93
rect 1936 47 1989 59
<< pdiff >>
rect 85 599 138 619
rect 85 565 93 599
rect 127 565 138 599
rect 85 505 138 565
rect 85 471 93 505
rect 127 471 138 505
rect 85 413 138 471
rect 85 379 93 413
rect 127 379 138 413
rect 85 367 138 379
rect 168 545 224 619
rect 168 511 179 545
rect 213 511 224 545
rect 168 477 224 511
rect 168 443 179 477
rect 213 443 224 477
rect 168 409 224 443
rect 168 375 179 409
rect 213 375 224 409
rect 168 367 224 375
rect 254 595 310 619
rect 254 561 265 595
rect 299 561 310 595
rect 254 518 310 561
rect 254 484 265 518
rect 299 484 310 518
rect 254 439 310 484
rect 254 405 265 439
rect 299 405 310 439
rect 254 367 310 405
rect 340 545 396 619
rect 340 511 351 545
rect 385 511 396 545
rect 340 477 396 511
rect 340 443 351 477
rect 385 443 396 477
rect 340 409 396 443
rect 340 375 351 409
rect 385 375 396 409
rect 340 367 396 375
rect 426 599 479 619
rect 426 565 437 599
rect 471 565 479 599
rect 426 518 479 565
rect 426 484 437 518
rect 471 484 479 518
rect 426 439 479 484
rect 426 405 437 439
rect 471 405 479 439
rect 426 367 479 405
rect 533 599 586 619
rect 533 565 541 599
rect 575 565 586 599
rect 533 495 586 565
rect 533 461 541 495
rect 575 461 586 495
rect 533 367 586 461
rect 616 504 672 619
rect 616 470 627 504
rect 661 470 672 504
rect 616 409 672 470
rect 616 375 627 409
rect 661 375 672 409
rect 616 367 672 375
rect 702 599 758 619
rect 702 565 713 599
rect 747 565 758 599
rect 702 367 758 565
rect 788 504 844 619
rect 788 470 799 504
rect 833 470 844 504
rect 788 367 844 470
rect 874 599 930 619
rect 874 565 885 599
rect 919 565 930 599
rect 874 367 930 565
rect 960 504 1016 619
rect 960 470 971 504
rect 1005 470 1016 504
rect 960 367 1016 470
rect 1046 599 1102 619
rect 1046 565 1057 599
rect 1091 565 1102 599
rect 1046 367 1102 565
rect 1132 504 1188 619
rect 1132 470 1143 504
rect 1177 470 1188 504
rect 1132 367 1188 470
rect 1218 599 1298 619
rect 1218 565 1241 599
rect 1275 565 1298 599
rect 1218 519 1298 565
rect 1218 485 1241 519
rect 1275 485 1298 519
rect 1218 447 1298 485
rect 1218 413 1253 447
rect 1287 413 1298 447
rect 1218 367 1298 413
rect 1328 607 1390 619
rect 1328 573 1341 607
rect 1375 573 1390 607
rect 1328 497 1390 573
rect 1328 463 1341 497
rect 1375 463 1390 497
rect 1328 367 1390 463
rect 1420 599 1476 619
rect 1420 565 1431 599
rect 1465 565 1476 599
rect 1420 512 1476 565
rect 1420 478 1431 512
rect 1465 478 1476 512
rect 1420 425 1476 478
rect 1420 391 1431 425
rect 1465 391 1476 425
rect 1420 367 1476 391
rect 1506 607 1562 619
rect 1506 573 1517 607
rect 1551 573 1562 607
rect 1506 497 1562 573
rect 1506 463 1517 497
rect 1551 463 1562 497
rect 1506 367 1562 463
rect 1592 599 1648 619
rect 1592 565 1603 599
rect 1637 565 1648 599
rect 1592 512 1648 565
rect 1592 478 1603 512
rect 1637 478 1648 512
rect 1592 425 1648 478
rect 1592 391 1603 425
rect 1637 391 1648 425
rect 1592 367 1648 391
rect 1678 607 1734 619
rect 1678 573 1689 607
rect 1723 573 1734 607
rect 1678 497 1734 573
rect 1678 463 1689 497
rect 1723 463 1734 497
rect 1678 367 1734 463
rect 1764 599 1820 619
rect 1764 565 1775 599
rect 1809 565 1820 599
rect 1764 505 1820 565
rect 1764 471 1775 505
rect 1809 471 1820 505
rect 1764 413 1820 471
rect 1764 379 1775 413
rect 1809 379 1820 413
rect 1764 367 1820 379
rect 1850 607 1906 619
rect 1850 573 1861 607
rect 1895 573 1906 607
rect 1850 512 1906 573
rect 1850 478 1861 512
rect 1895 478 1906 512
rect 1850 423 1906 478
rect 1850 389 1861 423
rect 1895 389 1906 423
rect 1850 367 1906 389
rect 1936 599 1989 619
rect 1936 565 1947 599
rect 1981 565 1989 599
rect 1936 505 1989 565
rect 1936 471 1947 505
rect 1981 471 1989 505
rect 1936 413 1989 471
rect 1936 379 1947 413
rect 1981 379 1989 413
rect 1936 367 1989 379
<< ndiffc >>
rect 127 169 161 203
rect 127 59 161 93
rect 213 158 247 192
rect 213 67 247 101
rect 299 98 333 132
rect 385 158 419 192
rect 385 67 419 101
rect 471 98 505 132
rect 557 117 591 151
rect 643 59 677 93
rect 729 67 763 101
rect 871 168 905 202
rect 957 67 991 101
rect 1043 168 1077 202
rect 1157 67 1191 101
rect 1243 96 1277 130
rect 1345 59 1379 93
rect 1431 156 1465 190
rect 1517 59 1551 93
rect 1603 156 1637 190
rect 1689 158 1723 192
rect 1689 67 1723 101
rect 1775 98 1809 132
rect 1861 158 1895 192
rect 1861 67 1895 101
rect 1947 169 1981 203
rect 1947 59 1981 93
<< pdiffc >>
rect 93 565 127 599
rect 93 471 127 505
rect 93 379 127 413
rect 179 511 213 545
rect 179 443 213 477
rect 179 375 213 409
rect 265 561 299 595
rect 265 484 299 518
rect 265 405 299 439
rect 351 511 385 545
rect 351 443 385 477
rect 351 375 385 409
rect 437 565 471 599
rect 437 484 471 518
rect 437 405 471 439
rect 541 565 575 599
rect 541 461 575 495
rect 627 470 661 504
rect 627 375 661 409
rect 713 565 747 599
rect 799 470 833 504
rect 885 565 919 599
rect 971 470 1005 504
rect 1057 565 1091 599
rect 1143 470 1177 504
rect 1241 565 1275 599
rect 1241 485 1275 519
rect 1253 413 1287 447
rect 1341 573 1375 607
rect 1341 463 1375 497
rect 1431 565 1465 599
rect 1431 478 1465 512
rect 1431 391 1465 425
rect 1517 573 1551 607
rect 1517 463 1551 497
rect 1603 565 1637 599
rect 1603 478 1637 512
rect 1603 391 1637 425
rect 1689 573 1723 607
rect 1689 463 1723 497
rect 1775 565 1809 599
rect 1775 471 1809 505
rect 1775 379 1809 413
rect 1861 573 1895 607
rect 1861 478 1895 512
rect 1861 389 1895 423
rect 1947 565 1981 599
rect 1947 471 1981 505
rect 1947 379 1981 413
<< poly >>
rect 138 619 168 645
rect 224 619 254 645
rect 310 619 340 645
rect 396 619 426 645
rect 586 619 616 645
rect 672 619 702 645
rect 758 619 788 645
rect 844 619 874 645
rect 930 619 960 645
rect 1016 619 1046 645
rect 1102 619 1132 645
rect 1188 619 1218 645
rect 1298 619 1328 645
rect 1390 619 1420 645
rect 1476 619 1506 645
rect 1562 619 1592 645
rect 1648 619 1678 645
rect 1734 619 1764 645
rect 1820 619 1850 645
rect 1906 619 1936 645
rect 138 303 168 367
rect 224 303 254 367
rect 310 303 340 367
rect 396 303 426 367
rect 586 335 616 367
rect 672 335 702 367
rect 758 335 788 367
rect 844 335 874 367
rect 930 335 960 367
rect 1016 335 1046 367
rect 1102 335 1132 367
rect 1188 335 1218 367
rect 1298 335 1328 367
rect 516 319 788 335
rect 45 287 460 303
rect 45 253 61 287
rect 95 253 129 287
rect 163 253 197 287
rect 231 253 265 287
rect 299 253 333 287
rect 367 253 401 287
rect 435 253 460 287
rect 45 237 460 253
rect 172 215 202 237
rect 258 215 288 237
rect 344 215 374 237
rect 430 215 460 237
rect 516 285 577 319
rect 611 285 645 319
rect 679 285 713 319
rect 747 285 788 319
rect 516 269 788 285
rect 830 319 1132 335
rect 830 285 846 319
rect 880 285 914 319
rect 948 285 982 319
rect 1016 285 1050 319
rect 1084 305 1132 319
rect 1174 319 1240 335
rect 1084 285 1118 305
rect 830 269 1118 285
rect 1174 285 1190 319
rect 1224 285 1240 319
rect 1174 269 1240 285
rect 1282 319 1348 335
rect 1282 285 1298 319
rect 1332 285 1348 319
rect 1282 269 1348 285
rect 1390 303 1420 367
rect 1476 303 1506 367
rect 1562 345 1592 367
rect 1648 345 1678 367
rect 1562 315 1678 345
rect 1562 303 1592 315
rect 1734 303 1764 367
rect 1820 303 1850 367
rect 1906 303 1936 367
rect 1390 287 1592 303
rect 516 215 546 269
rect 602 215 632 269
rect 688 215 718 269
rect 830 215 860 269
rect 916 215 946 269
rect 1002 215 1032 269
rect 1088 215 1118 269
rect 1202 215 1232 269
rect 1304 215 1334 269
rect 1390 253 1406 287
rect 1440 253 1474 287
rect 1508 253 1542 287
rect 1576 267 1592 287
rect 1720 287 1990 303
rect 1576 253 1678 267
rect 1390 237 1678 253
rect 1720 253 1736 287
rect 1770 253 1804 287
rect 1838 253 1872 287
rect 1906 253 1940 287
rect 1974 253 1990 287
rect 1720 237 1990 253
rect 1390 215 1420 237
rect 1476 215 1506 237
rect 1562 215 1592 237
rect 1648 215 1678 237
rect 1734 215 1764 237
rect 1820 215 1850 237
rect 1906 215 1936 237
rect 172 21 202 47
rect 258 21 288 47
rect 344 21 374 47
rect 430 21 460 47
rect 516 21 546 47
rect 602 21 632 47
rect 688 21 718 47
rect 830 21 860 47
rect 916 21 946 47
rect 1002 21 1032 47
rect 1088 21 1118 47
rect 1202 21 1232 47
rect 1304 21 1334 47
rect 1390 21 1420 47
rect 1476 21 1506 47
rect 1562 21 1592 47
rect 1648 21 1678 47
rect 1734 21 1764 47
rect 1820 21 1850 47
rect 1906 21 1936 47
<< polycont >>
rect 61 253 95 287
rect 129 253 163 287
rect 197 253 231 287
rect 265 253 299 287
rect 333 253 367 287
rect 401 253 435 287
rect 577 285 611 319
rect 645 285 679 319
rect 713 285 747 319
rect 846 285 880 319
rect 914 285 948 319
rect 982 285 1016 319
rect 1050 285 1084 319
rect 1190 285 1224 319
rect 1298 285 1332 319
rect 1406 253 1440 287
rect 1474 253 1508 287
rect 1542 253 1576 287
rect 1736 253 1770 287
rect 1804 253 1838 287
rect 1872 253 1906 287
rect 1940 253 1974 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 77 599 487 615
rect 77 565 93 599
rect 127 595 437 599
rect 127 581 265 595
rect 127 565 129 581
rect 77 505 129 565
rect 263 561 265 581
rect 299 581 437 595
rect 299 561 301 581
rect 77 471 93 505
rect 127 471 129 505
rect 77 413 129 471
rect 77 379 93 413
rect 127 379 129 413
rect 77 363 129 379
rect 163 545 229 547
rect 163 511 179 545
rect 213 511 229 545
rect 163 477 229 511
rect 163 443 179 477
rect 213 443 229 477
rect 163 409 229 443
rect 163 375 179 409
rect 213 375 229 409
rect 263 518 301 561
rect 435 565 437 581
rect 471 565 487 599
rect 263 484 265 518
rect 299 484 301 518
rect 263 439 301 484
rect 263 405 265 439
rect 299 405 301 439
rect 263 389 301 405
rect 335 545 401 547
rect 335 511 351 545
rect 385 511 401 545
rect 335 477 401 511
rect 335 443 351 477
rect 385 443 401 477
rect 335 409 401 443
rect 163 355 229 375
rect 335 375 351 409
rect 385 375 401 409
rect 435 518 487 565
rect 435 484 437 518
rect 471 484 487 518
rect 435 439 487 484
rect 525 599 1291 615
rect 525 565 541 599
rect 575 565 713 599
rect 747 565 885 599
rect 919 565 1057 599
rect 1091 565 1241 599
rect 1275 565 1291 599
rect 525 554 1291 565
rect 525 495 591 554
rect 525 461 541 495
rect 575 461 591 495
rect 525 457 591 461
rect 625 504 1193 520
rect 625 470 627 504
rect 661 470 799 504
rect 833 470 971 504
rect 1005 470 1143 504
rect 1177 470 1193 504
rect 435 405 437 439
rect 471 423 487 439
rect 625 454 1193 470
rect 1227 519 1291 554
rect 1227 485 1241 519
rect 1275 485 1291 519
rect 1227 454 1291 485
rect 1325 607 1391 649
rect 1325 573 1341 607
rect 1375 573 1391 607
rect 1325 497 1391 573
rect 1325 463 1341 497
rect 1375 463 1391 497
rect 1325 459 1391 463
rect 1427 599 1467 615
rect 1427 565 1431 599
rect 1465 565 1467 599
rect 1427 512 1467 565
rect 1427 478 1431 512
rect 1465 478 1467 512
rect 625 423 665 454
rect 471 409 665 423
rect 1251 447 1291 454
rect 471 405 627 409
rect 435 389 627 405
rect 335 355 401 375
rect 611 375 627 389
rect 661 375 665 409
rect 611 359 665 375
rect 729 386 1217 420
rect 1251 413 1253 447
rect 1287 425 1291 447
rect 1427 425 1467 478
rect 1501 607 1567 649
rect 1501 573 1517 607
rect 1551 573 1567 607
rect 1501 497 1567 573
rect 1501 463 1517 497
rect 1551 463 1567 497
rect 1501 459 1567 463
rect 1601 599 1639 615
rect 1601 565 1603 599
rect 1637 565 1639 599
rect 1601 512 1639 565
rect 1601 478 1603 512
rect 1637 478 1639 512
rect 1601 425 1639 478
rect 1673 607 1739 649
rect 1673 573 1689 607
rect 1723 573 1739 607
rect 1673 497 1739 573
rect 1673 463 1689 497
rect 1723 463 1739 497
rect 1673 459 1739 463
rect 1773 599 1811 615
rect 1773 565 1775 599
rect 1809 565 1811 599
rect 1773 505 1811 565
rect 1773 471 1775 505
rect 1809 471 1811 505
rect 1773 425 1811 471
rect 1287 413 1431 425
rect 1251 391 1431 413
rect 1465 391 1603 425
rect 1637 413 1811 425
rect 1637 391 1775 413
rect 163 321 527 355
rect 729 325 763 386
rect 17 253 61 287
rect 95 253 129 287
rect 163 253 197 287
rect 231 253 265 287
rect 299 253 333 287
rect 367 253 401 287
rect 435 253 453 287
rect 17 242 453 253
rect 487 251 527 321
rect 561 319 763 325
rect 561 285 577 319
rect 611 285 645 319
rect 679 285 713 319
rect 747 285 763 319
rect 797 319 1136 352
rect 797 285 846 319
rect 880 285 914 319
rect 948 285 982 319
rect 1016 285 1050 319
rect 1084 285 1136 319
rect 797 271 1136 285
rect 1170 335 1217 386
rect 1759 379 1775 391
rect 1809 379 1811 413
rect 1845 607 1911 649
rect 1845 573 1861 607
rect 1895 573 1911 607
rect 1845 512 1911 573
rect 1845 478 1861 512
rect 1895 478 1911 512
rect 1845 423 1911 478
rect 1845 389 1861 423
rect 1895 389 1911 423
rect 1945 599 1997 615
rect 1945 565 1947 599
rect 1981 565 1997 599
rect 1945 505 1997 565
rect 1945 471 1947 505
rect 1981 471 1997 505
rect 1945 413 1997 471
rect 1170 319 1240 335
rect 1170 285 1190 319
rect 1224 285 1240 319
rect 1170 269 1240 285
rect 1282 323 1697 357
rect 1282 319 1332 323
rect 1282 285 1298 319
rect 1649 287 1697 323
rect 1759 355 1811 379
rect 1945 379 1947 413
rect 1981 379 1997 413
rect 1945 355 1997 379
rect 1759 321 1997 355
rect 1282 269 1332 285
rect 1366 253 1406 287
rect 1440 253 1474 287
rect 1508 253 1542 287
rect 1576 253 1615 287
rect 487 237 763 251
rect 1366 240 1615 253
rect 1649 253 1736 287
rect 1770 253 1804 287
rect 1838 253 1872 287
rect 1906 253 1940 287
rect 1974 253 1999 287
rect 1649 242 1999 253
rect 487 208 1121 237
rect 111 203 177 208
rect 111 169 127 203
rect 161 169 177 203
rect 111 93 177 169
rect 111 59 127 93
rect 161 59 177 93
rect 111 17 177 59
rect 211 206 1121 208
rect 211 203 1651 206
rect 211 192 521 203
rect 211 158 213 192
rect 247 174 385 192
rect 247 158 249 174
rect 211 101 249 158
rect 383 158 385 174
rect 419 174 521 192
rect 797 202 1651 203
rect 419 158 421 174
rect 211 67 213 101
rect 247 67 249 101
rect 211 51 249 67
rect 283 132 349 140
rect 283 98 299 132
rect 333 98 349 132
rect 283 17 349 98
rect 383 101 421 158
rect 555 151 763 169
rect 797 168 871 202
rect 905 168 1043 202
rect 1077 190 1651 202
rect 1077 172 1431 190
rect 1077 168 1193 172
rect 797 151 1193 168
rect 1415 156 1431 172
rect 1465 156 1603 190
rect 1637 156 1651 190
rect 383 67 385 101
rect 419 67 421 101
rect 383 51 421 67
rect 455 132 521 140
rect 455 98 471 132
rect 505 98 521 132
rect 555 117 557 151
rect 591 135 763 151
rect 1415 140 1651 156
rect 1685 192 1897 208
rect 1685 158 1689 192
rect 1723 174 1861 192
rect 1723 158 1725 174
rect 591 117 593 135
rect 555 101 593 117
rect 727 117 763 135
rect 1227 130 1293 138
rect 727 101 1191 117
rect 455 17 521 98
rect 627 93 693 101
rect 627 59 643 93
rect 677 59 693 93
rect 627 17 693 59
rect 727 67 729 101
rect 763 67 957 101
rect 991 67 1157 101
rect 727 51 1191 67
rect 1227 96 1243 130
rect 1277 96 1293 130
rect 1685 106 1725 158
rect 1859 158 1861 174
rect 1895 158 1897 192
rect 1227 17 1293 96
rect 1329 101 1725 106
rect 1329 93 1689 101
rect 1329 59 1345 93
rect 1379 59 1517 93
rect 1551 67 1689 93
rect 1723 67 1725 101
rect 1551 59 1725 67
rect 1329 51 1725 59
rect 1759 132 1825 140
rect 1759 98 1775 132
rect 1809 98 1825 132
rect 1759 17 1825 98
rect 1859 101 1897 158
rect 1859 67 1861 101
rect 1895 67 1897 101
rect 1859 51 1897 67
rect 1931 203 1997 208
rect 1931 169 1947 203
rect 1981 169 1997 203
rect 1931 93 1997 169
rect 1931 59 1947 93
rect 1981 59 1997 93
rect 1931 17 1997 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3977276
string GDS_START 3960696
<< end >>
