magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 753 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 356 47 386 215
rect 428 47 458 215
rect 558 47 588 215
rect 644 47 674 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 356 367 386 619
rect 464 367 494 619
rect 560 367 590 619
rect 644 367 674 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 204 166 215
rect 110 170 121 204
rect 155 170 166 204
rect 110 101 166 170
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 131 356 215
rect 196 121 311 131
rect 196 87 207 121
rect 241 97 311 121
rect 345 97 356 131
rect 241 87 356 97
rect 196 47 356 87
rect 386 47 428 215
rect 458 195 558 215
rect 458 161 489 195
rect 523 161 558 195
rect 458 101 558 161
rect 458 67 489 101
rect 523 67 558 101
rect 458 47 558 67
rect 588 129 644 215
rect 588 95 599 129
rect 633 95 644 129
rect 588 47 644 95
rect 674 189 727 215
rect 674 155 685 189
rect 719 155 727 189
rect 674 101 727 155
rect 674 67 685 101
rect 719 67 727 101
rect 674 47 727 67
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 510 80 573
rect 27 476 35 510
rect 69 476 80 510
rect 27 413 80 476
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 599 166 619
rect 110 565 121 599
rect 155 565 166 599
rect 110 501 166 565
rect 110 467 121 501
rect 155 467 166 501
rect 110 413 166 467
rect 110 379 121 413
rect 155 379 166 413
rect 110 367 166 379
rect 196 607 249 619
rect 196 573 207 607
rect 241 573 249 607
rect 196 533 249 573
rect 196 499 207 533
rect 241 499 249 533
rect 196 459 249 499
rect 196 425 207 459
rect 241 425 249 459
rect 196 367 249 425
rect 303 599 356 619
rect 303 565 311 599
rect 345 565 356 599
rect 303 520 356 565
rect 303 486 311 520
rect 345 486 356 520
rect 303 443 356 486
rect 303 409 311 443
rect 345 409 356 443
rect 303 367 356 409
rect 386 607 464 619
rect 386 573 408 607
rect 442 573 464 607
rect 386 518 464 573
rect 386 484 408 518
rect 442 484 464 518
rect 386 367 464 484
rect 494 597 560 619
rect 494 563 508 597
rect 542 563 560 597
rect 494 518 560 563
rect 494 484 508 518
rect 542 484 560 518
rect 494 443 560 484
rect 494 409 508 443
rect 542 409 560 443
rect 494 367 560 409
rect 590 367 644 619
rect 674 607 727 619
rect 674 573 685 607
rect 719 573 727 607
rect 674 507 727 573
rect 674 473 685 507
rect 719 473 727 507
rect 674 413 727 473
rect 674 379 685 413
rect 719 379 727 413
rect 674 367 727 379
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 170 155 204
rect 121 67 155 101
rect 207 87 241 121
rect 311 97 345 131
rect 489 161 523 195
rect 489 67 523 101
rect 599 95 633 129
rect 685 155 719 189
rect 685 67 719 101
<< pdiffc >>
rect 35 573 69 607
rect 35 476 69 510
rect 35 379 69 413
rect 121 565 155 599
rect 121 467 155 501
rect 121 379 155 413
rect 207 573 241 607
rect 207 499 241 533
rect 207 425 241 459
rect 311 565 345 599
rect 311 486 345 520
rect 311 409 345 443
rect 408 573 442 607
rect 408 484 442 518
rect 508 563 542 597
rect 508 484 542 518
rect 508 409 542 443
rect 685 573 719 607
rect 685 473 719 507
rect 685 379 719 413
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 356 619 386 645
rect 464 619 494 645
rect 560 619 590 645
rect 644 619 674 645
rect 80 335 110 367
rect 166 335 196 367
rect 80 319 254 335
rect 80 285 204 319
rect 238 285 254 319
rect 356 305 386 367
rect 80 269 254 285
rect 303 289 386 305
rect 464 303 494 367
rect 560 303 590 367
rect 644 303 674 367
rect 80 215 110 269
rect 166 215 196 269
rect 303 255 319 289
rect 353 255 386 289
rect 303 239 386 255
rect 356 215 386 239
rect 428 287 494 303
rect 428 253 444 287
rect 478 253 494 287
rect 428 237 494 253
rect 536 287 602 303
rect 536 253 552 287
rect 586 253 602 287
rect 536 237 602 253
rect 644 287 743 303
rect 644 253 693 287
rect 727 253 743 287
rect 644 237 743 253
rect 428 215 458 237
rect 558 215 588 237
rect 644 215 674 237
rect 80 21 110 47
rect 166 21 196 47
rect 356 21 386 47
rect 428 21 458 47
rect 558 21 588 47
rect 644 21 674 47
<< polycont >>
rect 204 285 238 319
rect 319 255 353 289
rect 444 253 478 287
rect 552 253 586 287
rect 693 253 727 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 607 77 649
rect 19 573 35 607
rect 69 573 77 607
rect 19 510 77 573
rect 19 476 35 510
rect 69 476 77 510
rect 19 413 77 476
rect 19 379 35 413
rect 69 379 77 413
rect 19 363 77 379
rect 111 599 165 615
rect 111 565 121 599
rect 155 565 165 599
rect 111 501 165 565
rect 111 467 121 501
rect 155 467 165 501
rect 111 413 165 467
rect 111 379 121 413
rect 155 379 165 413
rect 200 607 257 649
rect 200 573 207 607
rect 241 573 257 607
rect 200 533 257 573
rect 200 499 207 533
rect 241 499 257 533
rect 200 459 257 499
rect 200 425 207 459
rect 241 425 257 459
rect 200 409 257 425
rect 295 599 358 615
rect 295 565 311 599
rect 345 565 358 599
rect 295 520 358 565
rect 295 486 311 520
rect 345 486 358 520
rect 295 445 358 486
rect 392 607 458 649
rect 392 573 408 607
rect 442 573 458 607
rect 392 518 458 573
rect 392 484 408 518
rect 442 484 458 518
rect 392 479 458 484
rect 492 597 558 613
rect 492 563 508 597
rect 542 563 558 597
rect 492 518 558 563
rect 492 484 508 518
rect 542 484 558 518
rect 492 445 558 484
rect 295 443 558 445
rect 295 409 311 443
rect 345 409 508 443
rect 542 409 558 443
rect 669 607 735 615
rect 669 573 685 607
rect 719 573 735 607
rect 669 507 735 573
rect 669 473 685 507
rect 719 473 735 507
rect 669 413 735 473
rect 19 203 77 219
rect 19 169 35 203
rect 69 169 77 203
rect 19 93 77 169
rect 19 59 35 93
rect 69 59 77 93
rect 19 17 77 59
rect 111 204 165 379
rect 669 379 685 413
rect 719 379 735 413
rect 669 375 735 379
rect 249 339 735 375
rect 249 335 283 339
rect 200 319 283 335
rect 200 285 204 319
rect 238 285 283 319
rect 200 269 283 285
rect 111 170 121 204
rect 155 170 165 204
rect 249 205 283 269
rect 317 289 369 305
rect 317 255 319 289
rect 353 255 369 289
rect 317 239 369 255
rect 403 287 494 303
rect 403 253 444 287
rect 478 253 494 287
rect 403 239 494 253
rect 536 287 643 303
rect 536 253 552 287
rect 586 253 643 287
rect 536 239 643 253
rect 677 287 751 303
rect 677 253 693 287
rect 727 253 751 287
rect 677 239 751 253
rect 249 195 735 205
rect 249 171 489 195
rect 111 101 165 170
rect 473 161 489 171
rect 523 189 735 195
rect 523 171 685 189
rect 523 161 539 171
rect 111 67 121 101
rect 155 67 165 101
rect 111 51 165 67
rect 199 131 361 137
rect 199 121 311 131
rect 199 87 207 121
rect 241 97 311 121
rect 345 97 361 131
rect 241 87 361 97
rect 199 17 361 87
rect 473 101 539 161
rect 683 155 685 171
rect 719 155 735 189
rect 473 67 489 101
rect 523 67 539 101
rect 473 51 539 67
rect 583 129 649 137
rect 583 95 599 129
rect 633 95 649 129
rect 583 17 649 95
rect 683 101 735 155
rect 683 67 685 101
rect 719 67 735 101
rect 683 51 735 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1961834
string GDS_START 1954194
<< end >>
