magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 5042 1975
<< nwell >>
rect -38 331 3782 704
rect 449 313 805 331
<< pwell >>
rect 476 229 977 249
rect 1 183 977 229
rect 1404 235 1911 279
rect 1404 229 2327 235
rect 2531 229 2639 275
rect 1404 207 2639 229
rect 1223 183 2639 207
rect 1 49 2639 183
rect 2920 182 3030 191
rect 3552 182 3743 241
rect 2920 49 3743 182
rect 0 0 3744 49
<< scnmos >>
rect 81 119 111 203
rect 159 119 189 203
rect 245 119 275 203
rect 339 119 369 203
rect 559 139 589 223
rect 659 139 689 223
rect 857 139 887 223
rect 966 73 996 157
rect 1068 47 1098 131
rect 1306 97 1336 181
rect 1385 97 1415 181
rect 1511 125 1541 253
rect 1626 125 1656 253
rect 1698 125 1728 253
rect 1900 125 1930 209
rect 1972 125 2002 209
rect 2044 125 2074 209
rect 2130 125 2160 209
rect 2216 125 2246 209
rect 2433 119 2463 203
rect 2505 119 2535 203
rect 3026 72 3056 156
rect 3104 72 3134 156
rect 3176 72 3206 156
rect 3262 72 3292 156
rect 3334 72 3364 156
rect 3526 47 3556 131
rect 3633 47 3663 215
<< scpmoshvt >>
rect 81 481 111 609
rect 183 481 213 609
rect 261 481 291 609
rect 347 481 377 609
rect 1016 535 1046 619
rect 1102 535 1132 619
rect 1180 535 1210 619
rect 1288 535 1318 619
rect 539 359 569 487
rect 685 359 715 487
rect 1397 451 1427 535
rect 1511 451 1541 619
rect 1682 451 1712 619
rect 1754 451 1784 619
rect 2470 401 2520 601
rect 2608 414 2658 614
rect 2706 414 2756 614
rect 2812 414 2862 614
rect 2916 414 2966 614
rect 3062 384 3092 512
rect 3148 384 3178 512
rect 3256 384 3306 584
rect 3523 403 3553 531
rect 3632 367 3662 619
<< ndiff >>
rect 27 178 81 203
rect 27 144 36 178
rect 70 144 81 178
rect 27 119 81 144
rect 111 119 159 203
rect 189 178 245 203
rect 189 144 200 178
rect 234 144 245 178
rect 189 119 245 144
rect 275 119 339 203
rect 369 178 434 203
rect 369 144 388 178
rect 422 144 434 178
rect 369 119 434 144
rect 502 185 559 223
rect 502 151 514 185
rect 548 151 559 185
rect 502 139 559 151
rect 589 185 659 223
rect 589 151 600 185
rect 634 151 659 185
rect 589 139 659 151
rect 689 198 746 223
rect 689 164 700 198
rect 734 164 746 198
rect 689 139 746 164
rect 800 206 857 223
rect 800 172 812 206
rect 846 172 857 206
rect 800 139 857 172
rect 887 198 951 223
rect 887 164 898 198
rect 932 164 951 198
rect 887 157 951 164
rect 887 139 966 157
rect 914 73 966 139
rect 996 131 1046 157
rect 1430 181 1511 253
rect 1249 169 1306 181
rect 1249 135 1261 169
rect 1295 135 1306 169
rect 996 73 1068 131
rect 1018 47 1068 73
rect 1098 97 1155 131
rect 1249 97 1306 135
rect 1336 97 1385 181
rect 1415 159 1511 181
rect 1415 125 1439 159
rect 1473 125 1511 159
rect 1541 237 1626 253
rect 1541 203 1581 237
rect 1615 203 1626 237
rect 1541 169 1626 203
rect 1541 135 1581 169
rect 1615 135 1626 169
rect 1541 125 1626 135
rect 1656 125 1698 253
rect 1728 245 1885 253
rect 1728 211 1789 245
rect 1823 211 1885 245
rect 1728 209 1885 211
rect 1728 125 1900 209
rect 1930 125 1972 209
rect 2002 125 2044 209
rect 2074 184 2130 209
rect 2074 150 2085 184
rect 2119 150 2130 184
rect 2074 125 2130 150
rect 2160 181 2216 209
rect 2160 147 2171 181
rect 2205 147 2216 181
rect 2160 125 2216 147
rect 2246 184 2301 209
rect 2557 237 2613 249
rect 2557 203 2569 237
rect 2603 203 2613 237
rect 2246 150 2257 184
rect 2291 150 2301 184
rect 2246 125 2301 150
rect 2355 170 2433 203
rect 2355 136 2365 170
rect 2399 136 2433 170
rect 1415 97 1489 125
rect 1098 63 1109 97
rect 1143 63 1155 97
rect 1098 47 1155 63
rect 2355 119 2433 136
rect 2463 119 2505 203
rect 2535 119 2613 203
rect 2946 156 3004 165
rect 2946 153 3026 156
rect 2946 119 2958 153
rect 2992 119 3026 153
rect 2946 72 3026 119
rect 3056 72 3104 156
rect 3134 72 3176 156
rect 3206 122 3262 156
rect 3206 88 3217 122
rect 3251 88 3262 122
rect 3206 72 3262 88
rect 3292 72 3334 156
rect 3364 131 3418 156
rect 3578 187 3633 215
rect 3578 153 3588 187
rect 3622 153 3633 187
rect 3578 131 3633 153
rect 3364 97 3375 131
rect 3409 97 3418 131
rect 3364 72 3418 97
rect 3472 106 3526 131
rect 3472 72 3481 106
rect 3515 72 3526 106
rect 3472 47 3526 72
rect 3556 93 3633 131
rect 3556 59 3588 93
rect 3622 59 3633 93
rect 3556 47 3633 59
rect 3663 203 3717 215
rect 3663 169 3674 203
rect 3708 169 3717 203
rect 3663 101 3717 169
rect 3663 67 3674 101
rect 3708 67 3717 101
rect 3663 47 3717 67
<< pdiff >>
rect 27 597 81 609
rect 27 563 36 597
rect 70 563 81 597
rect 27 527 81 563
rect 27 493 36 527
rect 70 493 81 527
rect 27 481 81 493
rect 111 597 183 609
rect 111 563 136 597
rect 170 563 183 597
rect 111 527 183 563
rect 111 493 136 527
rect 170 493 183 527
rect 111 481 183 493
rect 213 481 261 609
rect 291 537 347 609
rect 291 503 302 537
rect 336 503 347 537
rect 291 481 347 503
rect 377 580 431 609
rect 945 590 1016 619
rect 377 546 388 580
rect 422 546 431 580
rect 377 481 431 546
rect 591 563 643 575
rect 591 529 600 563
rect 634 529 643 563
rect 591 487 643 529
rect 945 556 957 590
rect 991 556 1016 590
rect 945 535 1016 556
rect 1046 590 1102 619
rect 1046 556 1057 590
rect 1091 556 1102 590
rect 1046 535 1102 556
rect 1132 535 1180 619
rect 1210 594 1288 619
rect 1210 560 1221 594
rect 1255 560 1288 594
rect 1210 535 1288 560
rect 1318 535 1382 619
rect 1454 607 1511 619
rect 1454 573 1466 607
rect 1500 573 1511 607
rect 1454 535 1511 573
rect 485 405 539 487
rect 485 371 494 405
rect 528 371 539 405
rect 485 359 539 371
rect 569 359 685 487
rect 715 405 769 487
rect 715 371 726 405
rect 760 371 769 405
rect 715 359 769 371
rect 1340 513 1397 535
rect 1340 479 1352 513
rect 1386 479 1397 513
rect 1340 451 1397 479
rect 1427 501 1511 535
rect 1427 467 1466 501
rect 1500 467 1511 501
rect 1427 451 1511 467
rect 1541 497 1682 619
rect 1541 463 1637 497
rect 1671 463 1682 497
rect 1541 451 1682 463
rect 1712 451 1754 619
rect 1784 590 1841 619
rect 1784 556 1795 590
rect 1829 556 1841 590
rect 1784 497 1841 556
rect 2535 615 2593 627
rect 2535 601 2547 615
rect 1784 463 1795 497
rect 1829 463 1841 497
rect 1784 451 1841 463
rect 2299 447 2470 601
rect 2299 413 2311 447
rect 2345 413 2470 447
rect 2299 401 2470 413
rect 2520 581 2547 601
rect 2581 614 2593 615
rect 2581 581 2608 614
rect 2520 414 2608 581
rect 2658 414 2706 614
rect 2756 525 2812 614
rect 2756 491 2767 525
rect 2801 491 2812 525
rect 2756 414 2812 491
rect 2862 414 2916 614
rect 2966 590 3040 614
rect 2966 556 2997 590
rect 3031 556 3040 590
rect 3575 607 3632 619
rect 2966 512 3040 556
rect 3200 569 3256 584
rect 3200 535 3211 569
rect 3245 535 3256 569
rect 3200 512 3256 535
rect 2966 414 3062 512
rect 2520 401 2570 414
rect 2988 384 3062 414
rect 3092 430 3148 512
rect 3092 396 3103 430
rect 3137 396 3148 430
rect 3092 384 3148 396
rect 3178 384 3256 512
rect 3306 430 3363 584
rect 3575 573 3587 607
rect 3621 573 3632 607
rect 3575 531 3632 573
rect 3306 396 3317 430
rect 3351 396 3363 430
rect 3466 519 3523 531
rect 3466 485 3478 519
rect 3512 485 3523 519
rect 3466 449 3523 485
rect 3466 415 3478 449
rect 3512 415 3523 449
rect 3466 403 3523 415
rect 3553 510 3632 531
rect 3553 476 3587 510
rect 3621 476 3632 510
rect 3553 413 3632 476
rect 3553 403 3587 413
rect 3306 384 3363 396
rect 3575 379 3587 403
rect 3621 379 3632 413
rect 3575 367 3632 379
rect 3662 599 3717 619
rect 3662 565 3673 599
rect 3707 565 3717 599
rect 3662 506 3717 565
rect 3662 472 3673 506
rect 3707 472 3717 506
rect 3662 413 3717 472
rect 3662 379 3673 413
rect 3707 379 3717 413
rect 3662 367 3717 379
<< ndiffc >>
rect 36 144 70 178
rect 200 144 234 178
rect 388 144 422 178
rect 514 151 548 185
rect 600 151 634 185
rect 700 164 734 198
rect 812 172 846 206
rect 898 164 932 198
rect 1261 135 1295 169
rect 1439 125 1473 159
rect 1581 203 1615 237
rect 1581 135 1615 169
rect 1789 211 1823 245
rect 2085 150 2119 184
rect 2171 147 2205 181
rect 2569 203 2603 237
rect 2257 150 2291 184
rect 2365 136 2399 170
rect 1109 63 1143 97
rect 2958 119 2992 153
rect 3217 88 3251 122
rect 3588 153 3622 187
rect 3375 97 3409 131
rect 3481 72 3515 106
rect 3588 59 3622 93
rect 3674 169 3708 203
rect 3674 67 3708 101
<< pdiffc >>
rect 36 563 70 597
rect 36 493 70 527
rect 136 563 170 597
rect 136 493 170 527
rect 302 503 336 537
rect 388 546 422 580
rect 600 529 634 563
rect 957 556 991 590
rect 1057 556 1091 590
rect 1221 560 1255 594
rect 1466 573 1500 607
rect 494 371 528 405
rect 726 371 760 405
rect 1352 479 1386 513
rect 1466 467 1500 501
rect 1637 463 1671 497
rect 1795 556 1829 590
rect 1795 463 1829 497
rect 2311 413 2345 447
rect 2547 581 2581 615
rect 2767 491 2801 525
rect 2997 556 3031 590
rect 3211 535 3245 569
rect 3103 396 3137 430
rect 3587 573 3621 607
rect 3317 396 3351 430
rect 3478 485 3512 519
rect 3478 415 3512 449
rect 3587 476 3621 510
rect 3587 379 3621 413
rect 3673 565 3707 599
rect 3673 472 3707 506
rect 3673 379 3707 413
<< poly >>
rect 81 609 111 635
rect 183 609 213 635
rect 261 609 291 635
rect 347 609 377 635
rect 1016 619 1046 645
rect 1102 619 1132 645
rect 1180 619 1210 645
rect 1288 619 1318 645
rect 1511 619 1541 645
rect 1682 619 1712 645
rect 1754 619 1784 645
rect 539 487 569 513
rect 685 487 715 585
rect 1397 535 1427 561
rect 81 375 111 481
rect 183 447 213 481
rect 45 359 111 375
rect 45 325 61 359
rect 95 325 111 359
rect 45 291 111 325
rect 45 257 61 291
rect 95 257 111 291
rect 45 241 111 257
rect 81 203 111 241
rect 153 417 213 447
rect 153 255 183 417
rect 261 375 291 481
rect 347 395 377 481
rect 225 359 291 375
rect 225 325 241 359
rect 275 325 291 359
rect 225 309 291 325
rect 339 379 453 395
rect 339 345 403 379
rect 437 345 453 379
rect 1016 479 1046 535
rect 801 463 1046 479
rect 801 429 817 463
rect 851 449 1046 463
rect 851 429 867 449
rect 801 395 867 429
rect 801 361 817 395
rect 851 361 867 395
rect 339 311 453 345
rect 153 225 189 255
rect 159 203 189 225
rect 245 203 275 309
rect 339 277 403 311
rect 437 277 453 311
rect 339 261 453 277
rect 539 311 569 359
rect 539 295 611 311
rect 539 261 561 295
rect 595 261 611 295
rect 685 275 715 359
rect 801 345 867 361
rect 1102 291 1132 535
rect 1180 503 1210 535
rect 1180 487 1246 503
rect 1180 453 1196 487
rect 1230 453 1246 487
rect 1180 437 1246 453
rect 1090 275 1156 291
rect 339 203 369 261
rect 539 245 611 261
rect 659 245 1106 275
rect 559 223 589 245
rect 659 223 689 245
rect 857 223 887 245
rect 1090 241 1106 245
rect 1140 241 1156 275
rect 1216 269 1246 437
rect 1288 419 1318 535
rect 2201 599 2275 615
rect 2470 601 2520 627
rect 2201 565 2217 599
rect 2251 565 2275 599
rect 2201 549 2275 565
rect 1288 403 1354 419
rect 1288 369 1304 403
rect 1338 369 1354 403
rect 1288 353 1354 369
rect 1090 225 1156 241
rect 1198 253 1264 269
rect 1198 219 1214 253
rect 1248 219 1264 253
rect 1198 203 1264 219
rect 1198 183 1228 203
rect 966 157 996 183
rect 81 93 111 119
rect 159 51 189 119
rect 245 93 275 119
rect 339 93 369 119
rect 559 51 589 139
rect 659 113 689 139
rect 159 21 589 51
rect 737 101 803 117
rect 857 113 887 139
rect 737 67 753 101
rect 787 67 803 101
rect 1068 153 1228 183
rect 1306 181 1336 353
rect 1397 298 1427 451
rect 1511 419 1541 451
rect 1469 403 1541 419
rect 1469 369 1485 403
rect 1519 369 1541 403
rect 1682 429 1712 451
rect 1754 429 1784 451
rect 1682 413 2083 429
rect 1682 399 2033 413
rect 1469 321 1541 369
rect 1385 268 1427 298
rect 1385 181 1415 268
rect 1511 253 1541 321
rect 1626 332 1762 348
rect 1626 298 1712 332
rect 1746 298 1762 332
rect 1626 282 1762 298
rect 1626 253 1656 282
rect 1698 253 1728 282
rect 1068 131 1098 153
rect 737 51 803 67
rect 966 51 996 73
rect 737 21 996 51
rect 1900 209 1930 399
rect 2017 379 2033 399
rect 2067 379 2083 413
rect 2017 363 2083 379
rect 2131 427 2197 443
rect 2131 393 2147 427
rect 2181 393 2197 427
rect 2131 377 2197 393
rect 2245 379 2275 549
rect 2608 614 2658 640
rect 2706 614 2756 640
rect 2812 614 2862 640
rect 2916 614 2966 640
rect 3632 619 3662 645
rect 3256 584 3306 610
rect 3062 512 3092 538
rect 3148 512 3178 538
rect 2470 379 2520 401
rect 2131 315 2161 377
rect 2245 349 2535 379
rect 1972 285 2161 315
rect 1972 209 2002 285
rect 2044 209 2074 285
rect 2325 275 2391 291
rect 2325 261 2341 275
rect 2216 241 2341 261
rect 2375 241 2391 275
rect 2130 209 2160 235
rect 2216 231 2391 241
rect 2216 209 2246 231
rect 2325 225 2391 231
rect 2433 203 2463 349
rect 2505 203 2535 349
rect 2608 274 2658 414
rect 2706 384 2756 414
rect 2700 366 2766 384
rect 2812 382 2862 414
rect 2916 388 2966 414
rect 2700 332 2716 366
rect 2750 332 2766 366
rect 2700 316 2766 332
rect 2808 366 2874 382
rect 2808 332 2824 366
rect 2858 332 2874 366
rect 2808 316 2874 332
rect 2608 264 2694 274
rect 2628 244 2694 264
rect 1511 99 1541 125
rect 1626 99 1656 125
rect 1698 99 1728 125
rect 1900 99 1930 125
rect 1972 99 2002 125
rect 2044 99 2074 125
rect 1306 71 1336 97
rect 1385 51 1415 97
rect 2130 51 2160 125
rect 2216 99 2246 125
rect 2664 159 2694 244
rect 2736 268 2766 316
rect 2916 274 2951 388
rect 3523 531 3553 557
rect 3062 335 3092 384
rect 2736 238 2843 268
rect 2664 143 2771 159
rect 2433 93 2463 119
rect 2505 93 2535 119
rect 2664 109 2721 143
rect 2755 109 2771 143
rect 2664 93 2771 109
rect 2813 51 2843 238
rect 2885 258 2951 274
rect 2993 319 3092 335
rect 2993 285 3009 319
rect 3043 285 3092 319
rect 3148 310 3178 384
rect 3256 358 3306 384
rect 3523 381 3553 403
rect 3437 365 3553 381
rect 3276 310 3306 358
rect 2993 269 3092 285
rect 3134 294 3306 310
rect 3401 351 3553 365
rect 3401 349 3467 351
rect 3401 315 3417 349
rect 3451 315 3467 349
rect 3401 299 3467 315
rect 3632 303 3662 367
rect 2885 224 2901 258
rect 2935 224 2951 258
rect 2885 208 2951 224
rect 3026 156 3056 269
rect 3134 260 3202 294
rect 3236 260 3306 294
rect 3134 251 3306 260
rect 3134 221 3364 251
rect 3104 191 3206 221
rect 3104 156 3134 191
rect 3176 156 3206 191
rect 3262 156 3292 221
rect 3334 156 3364 221
rect 3437 189 3467 299
rect 3586 287 3663 303
rect 3586 253 3602 287
rect 3636 253 3663 287
rect 3586 237 3663 253
rect 3633 215 3663 237
rect 3437 159 3556 189
rect 3526 131 3556 159
rect 1068 21 1098 47
rect 1385 21 2843 51
rect 3026 46 3056 72
rect 3104 46 3134 72
rect 3176 46 3206 72
rect 3262 46 3292 72
rect 3334 46 3364 72
rect 3526 21 3556 47
rect 3633 21 3663 47
<< polycont >>
rect 61 325 95 359
rect 61 257 95 291
rect 241 325 275 359
rect 403 345 437 379
rect 817 429 851 463
rect 817 361 851 395
rect 403 277 437 311
rect 561 261 595 295
rect 1196 453 1230 487
rect 1106 241 1140 275
rect 2217 565 2251 599
rect 1304 369 1338 403
rect 1214 219 1248 253
rect 753 67 787 101
rect 1485 369 1519 403
rect 1712 298 1746 332
rect 2033 379 2067 413
rect 2147 393 2181 427
rect 2341 241 2375 275
rect 2716 332 2750 366
rect 2824 332 2858 366
rect 2721 109 2755 143
rect 3009 285 3043 319
rect 3417 315 3451 349
rect 2901 224 2935 258
rect 3202 260 3236 294
rect 3602 253 3636 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3744 683
rect 20 597 86 613
rect 20 563 36 597
rect 70 563 86 597
rect 20 527 86 563
rect 20 493 36 527
rect 70 493 86 527
rect 20 443 86 493
rect 120 597 170 649
rect 120 563 136 597
rect 120 527 170 563
rect 120 493 136 527
rect 120 477 170 493
rect 204 581 438 615
rect 204 443 238 581
rect 388 580 438 581
rect 286 537 354 547
rect 286 503 302 537
rect 336 503 354 537
rect 422 546 438 580
rect 388 513 438 546
rect 584 563 650 649
rect 920 590 1007 615
rect 920 565 957 590
rect 584 529 600 563
rect 634 529 650 563
rect 584 513 650 529
rect 733 556 957 565
rect 991 556 1007 590
rect 733 531 1007 556
rect 1041 590 1107 615
rect 1041 556 1057 590
rect 1091 556 1107 590
rect 286 479 354 503
rect 733 479 767 531
rect 286 445 767 479
rect 801 463 852 479
rect 20 409 238 443
rect 25 359 167 375
rect 25 325 61 359
rect 95 325 167 359
rect 25 291 167 325
rect 217 359 286 375
rect 217 325 241 359
rect 275 325 286 359
rect 217 309 286 325
rect 25 257 61 291
rect 95 257 167 291
rect 25 241 167 257
rect 320 207 354 445
rect 801 429 817 463
rect 851 429 852 463
rect 801 411 852 429
rect 388 405 544 411
rect 388 379 494 405
rect 388 345 403 379
rect 437 371 494 379
rect 528 371 544 405
rect 437 345 544 371
rect 684 405 852 411
rect 684 371 726 405
rect 760 395 852 405
rect 760 371 817 395
rect 684 361 817 371
rect 851 361 852 395
rect 684 345 852 361
rect 388 311 511 345
rect 388 277 403 311
rect 437 277 511 311
rect 388 261 511 277
rect 20 178 86 207
rect 20 144 36 178
rect 70 144 86 178
rect 20 17 86 144
rect 184 178 354 207
rect 184 144 200 178
rect 234 173 354 178
rect 388 178 438 207
rect 234 144 250 173
rect 184 115 250 144
rect 422 144 438 178
rect 388 17 438 144
rect 477 202 511 261
rect 545 295 647 311
rect 545 261 561 295
rect 595 261 647 295
rect 545 236 647 261
rect 477 185 548 202
rect 477 151 514 185
rect 477 135 548 151
rect 584 185 650 202
rect 584 151 600 185
rect 634 151 650 185
rect 584 17 650 151
rect 684 198 750 345
rect 886 311 920 531
rect 1041 415 1107 556
rect 1205 594 1271 649
rect 1205 560 1221 594
rect 1255 560 1271 594
rect 1205 531 1271 560
rect 1450 607 1516 649
rect 1450 573 1466 607
rect 1500 573 1516 607
rect 1551 581 1739 615
rect 1336 513 1402 539
rect 1336 497 1352 513
rect 1180 487 1352 497
rect 1180 453 1196 487
rect 1230 479 1352 487
rect 1386 479 1402 513
rect 1230 453 1402 479
rect 1450 501 1516 573
rect 1450 467 1466 501
rect 1500 467 1516 501
rect 1450 453 1516 467
rect 1180 449 1246 453
rect 1288 415 1535 419
rect 684 164 700 198
rect 734 164 750 198
rect 684 117 750 164
rect 796 277 920 311
rect 954 403 1535 415
rect 954 381 1304 403
rect 796 206 846 277
rect 954 227 988 381
rect 1288 369 1304 381
rect 1338 369 1485 403
rect 1519 369 1535 403
rect 1288 362 1535 369
rect 796 172 812 206
rect 796 151 846 172
rect 882 198 988 227
rect 882 164 898 198
rect 932 164 988 198
rect 882 135 988 164
rect 1022 328 1224 343
rect 1569 328 1603 581
rect 1022 309 1603 328
rect 684 101 803 117
rect 684 67 753 101
rect 787 85 803 101
rect 1022 85 1056 309
rect 1190 294 1603 309
rect 1637 497 1671 513
rect 1090 241 1106 275
rect 1140 241 1156 275
rect 1090 169 1156 241
rect 1198 253 1311 260
rect 1198 219 1214 253
rect 1248 219 1311 253
rect 1198 203 1311 219
rect 1261 169 1311 203
rect 1090 135 1227 169
rect 787 67 1056 85
rect 684 51 1056 67
rect 1093 97 1159 101
rect 1093 63 1109 97
rect 1143 63 1159 97
rect 1093 17 1159 63
rect 1193 85 1227 135
rect 1295 135 1311 169
rect 1261 119 1311 135
rect 1345 226 1541 260
rect 1637 253 1671 463
rect 1345 85 1379 226
rect 1193 51 1379 85
rect 1423 159 1473 192
rect 1423 125 1439 159
rect 1423 17 1473 125
rect 1507 85 1541 226
rect 1575 237 1671 253
rect 1575 203 1581 237
rect 1615 219 1671 237
rect 1705 348 1739 581
rect 1788 599 2497 615
rect 1788 590 2217 599
rect 1788 556 1795 590
rect 1829 565 2217 590
rect 2251 565 2497 599
rect 2531 581 2547 615
rect 2581 590 3047 615
rect 2581 581 2997 590
rect 3031 581 3047 590
rect 3571 607 3637 649
rect 1829 556 2497 565
rect 1788 549 2497 556
rect 1779 497 1829 549
rect 2463 547 2497 549
rect 2981 556 2997 581
rect 2981 547 3007 556
rect 3041 547 3047 581
rect 2463 525 2826 547
rect 2981 532 3047 547
rect 3193 581 3261 588
rect 3193 547 3199 581
rect 3233 569 3261 581
rect 3193 535 3211 547
rect 3245 535 3261 569
rect 3571 573 3587 607
rect 3621 573 3637 607
rect 3193 532 3261 535
rect 1779 463 1795 497
rect 1779 447 1829 463
rect 1863 481 2429 515
rect 2463 513 2767 525
rect 1705 332 1751 348
rect 1705 298 1712 332
rect 1746 298 1751 332
rect 1705 282 1751 298
rect 1615 203 1629 219
rect 1575 169 1629 203
rect 1575 135 1581 169
rect 1615 135 1629 169
rect 1575 119 1629 135
rect 1705 153 1739 282
rect 1785 245 1819 447
rect 1863 427 1897 481
rect 2395 479 2429 481
rect 2760 491 2767 513
rect 2801 504 2826 525
rect 3478 519 3535 535
rect 2801 498 2919 504
rect 2801 491 3444 498
rect 1863 377 1907 427
rect 1773 211 1789 245
rect 1823 211 1839 245
rect 1773 187 1839 211
rect 1873 153 1907 377
rect 2033 413 2083 429
rect 2067 379 2083 413
rect 2033 343 2083 379
rect 2131 427 2197 443
rect 2131 393 2147 427
rect 2181 411 2197 427
rect 2295 413 2311 447
rect 2345 413 2361 447
rect 2395 445 2671 479
rect 2760 470 3444 491
rect 2885 464 3444 470
rect 2295 411 2361 413
rect 2637 436 2671 445
rect 2181 393 2603 411
rect 2637 402 2842 436
rect 2131 377 2603 393
rect 1705 119 1907 153
rect 2017 309 2535 343
rect 2017 85 2051 309
rect 2085 241 2291 275
rect 2085 184 2119 241
rect 2085 121 2119 150
rect 2155 181 2205 207
rect 2155 147 2171 181
rect 1507 51 2051 85
rect 2155 17 2205 147
rect 2241 184 2291 241
rect 2325 241 2341 275
rect 2375 241 2467 275
rect 2325 225 2467 241
rect 2241 150 2257 184
rect 2241 121 2291 150
rect 2349 170 2399 191
rect 2349 136 2365 170
rect 2349 17 2399 136
rect 2433 85 2467 225
rect 2501 153 2535 309
rect 2569 282 2603 377
rect 2808 382 2842 402
rect 2700 366 2766 368
rect 2700 332 2716 366
rect 2750 332 2766 366
rect 2700 316 2766 332
rect 2808 366 2874 382
rect 2808 332 2824 366
rect 2858 332 2874 366
rect 2808 316 2874 332
rect 2993 319 3047 430
rect 2993 285 3009 319
rect 3043 285 3047 319
rect 2569 258 2951 282
rect 2569 248 2901 258
rect 2569 237 2603 248
rect 2885 224 2901 248
rect 2935 224 2951 258
rect 2993 236 3047 285
rect 3081 396 3103 430
rect 3137 396 3153 430
rect 3081 380 3153 396
rect 2569 187 2603 203
rect 2637 180 2851 214
rect 2885 208 2951 224
rect 2637 153 2671 180
rect 2501 119 2671 153
rect 2817 169 2851 180
rect 3081 169 3115 380
rect 3187 294 3252 430
rect 3187 260 3202 294
rect 3236 260 3252 294
rect 3187 244 3252 260
rect 3291 396 3317 430
rect 3351 396 3367 430
rect 3291 210 3367 396
rect 3410 365 3444 464
rect 3512 485 3535 519
rect 3478 449 3535 485
rect 3512 415 3535 449
rect 3478 399 3535 415
rect 3401 349 3467 365
rect 3401 315 3417 349
rect 3451 315 3467 349
rect 3401 299 3467 315
rect 3501 303 3535 399
rect 3571 510 3637 573
rect 3571 476 3587 510
rect 3621 476 3637 510
rect 3571 413 3637 476
rect 3571 379 3587 413
rect 3621 379 3637 413
rect 3571 363 3637 379
rect 3673 599 3724 615
rect 3707 565 3724 599
rect 3673 506 3724 565
rect 3707 472 3724 506
rect 3673 413 3724 472
rect 3707 379 3724 413
rect 2817 153 3115 169
rect 2705 143 2771 146
rect 2705 109 2721 143
rect 2755 109 2771 143
rect 2817 119 2958 153
rect 2992 119 3115 153
rect 3149 176 3367 210
rect 2705 85 2771 109
rect 3149 85 3183 176
rect 3333 160 3367 176
rect 3501 287 3639 303
rect 3501 253 3602 287
rect 3636 253 3639 287
rect 3501 237 3639 253
rect 2433 51 3183 85
rect 3217 122 3267 142
rect 3333 131 3425 160
rect 3501 135 3535 237
rect 3673 203 3724 379
rect 3333 126 3375 131
rect 3251 88 3267 122
rect 3217 17 3267 88
rect 3359 97 3375 126
rect 3409 97 3425 131
rect 3359 84 3425 97
rect 3465 106 3535 135
rect 3465 72 3481 106
rect 3515 72 3535 106
rect 3465 59 3535 72
rect 3572 187 3638 203
rect 3572 153 3588 187
rect 3622 153 3638 187
rect 3572 93 3638 153
rect 3572 59 3588 93
rect 3622 59 3638 93
rect 3572 17 3638 59
rect 3673 169 3674 203
rect 3708 169 3724 203
rect 3673 101 3724 169
rect 3673 67 3674 101
rect 3708 67 3724 101
rect 3673 51 3724 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3007 556 3031 581
rect 3031 556 3041 581
rect 3007 547 3041 556
rect 3199 569 3233 581
rect 3199 547 3211 569
rect 3211 547 3233 569
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
<< metal1 >>
rect 0 683 3744 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3744 683
rect 0 617 3744 649
rect 14 581 3730 589
rect 14 547 3007 581
rect 3041 547 3199 581
rect 3233 547 3730 581
rect 14 535 3730 547
rect 0 17 3744 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
rect 0 -49 3744 -17
<< labels >>
flabel pwell s 0 0 3744 49 0 FreeSans 200 0 0 0 VNB
port 9 nsew ground bidirectional
flabel nwell s 0 617 3744 666 0 FreeSans 200 0 0 0 VPB
port 10 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srsdfstp_1
flabel comment s 1226 358 1226 358 0 FreeSans 200 90 0 0 no_jumper_check
flabel locali s 3679 242 3713 276 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 538 3713 572 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 464 3713 498 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 390 3713 424 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 316 3713 350 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 94 3713 128 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 3679 168 3713 202 0 FreeSans 200 0 0 0 Q
port 12 nsew signal output
flabel locali s 2719 316 2753 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3007 316 3041 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3199 316 3233 350 0 FreeSans 340 0 0 0 SLEEP_B
port 6 nsew signal input
flabel locali s 3199 390 3233 424 0 FreeSans 340 0 0 0 SLEEP_B
port 6 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel metal1 s 14 535 3730 589 0 FreeSans 340 0 0 0 KAPWR
port 7 nsew power bidirectional
flabel metal1 s 0 617 3744 666 0 FreeSans 200 0 0 0 VPWR
port 11 nsew power bidirectional
flabel metal1 s 0 0 3744 17 0 FreeSans 200 0 0 0 VGND
port 8 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3744 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2737552
string GDS_START 2712668
<< end >>
