magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 413 228 766 248
rect 1 49 766 228
rect 0 0 768 49
<< scpmos >>
rect 86 392 116 592
rect 170 392 200 592
rect 284 392 314 592
rect 535 368 565 536
rect 652 368 682 592
<< nmoslvt >>
rect 84 74 114 202
rect 198 74 228 202
rect 287 74 317 202
rect 539 112 569 222
rect 653 74 683 222
<< ndiff >>
rect 27 188 84 202
rect 27 154 39 188
rect 73 154 84 188
rect 27 120 84 154
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 122 198 202
rect 114 88 139 122
rect 173 88 198 122
rect 114 74 198 88
rect 228 188 287 202
rect 228 154 239 188
rect 273 154 287 188
rect 228 120 287 154
rect 228 86 239 120
rect 273 86 287 120
rect 228 74 287 86
rect 317 190 385 202
rect 317 156 339 190
rect 373 156 385 190
rect 317 120 385 156
rect 317 86 339 120
rect 373 86 385 120
rect 439 186 539 222
rect 439 152 494 186
rect 528 152 539 186
rect 439 112 539 152
rect 569 195 653 222
rect 569 161 594 195
rect 628 161 653 195
rect 569 116 653 161
rect 569 112 608 116
rect 317 74 385 86
rect 591 82 608 112
rect 642 82 653 116
rect 591 74 653 82
rect 683 210 740 222
rect 683 176 694 210
rect 728 176 740 210
rect 683 120 740 176
rect 683 86 694 120
rect 728 86 740 120
rect 683 74 740 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 512 86 546
rect 27 478 39 512
rect 73 478 86 512
rect 27 444 86 478
rect 27 410 39 444
rect 73 410 86 444
rect 27 392 86 410
rect 116 392 170 592
rect 200 580 284 592
rect 200 546 227 580
rect 261 546 284 580
rect 200 512 284 546
rect 200 478 227 512
rect 261 478 284 512
rect 200 444 284 478
rect 200 410 227 444
rect 261 410 284 444
rect 200 392 284 410
rect 314 573 373 592
rect 314 539 327 573
rect 361 539 373 573
rect 583 573 652 592
rect 314 392 373 539
rect 583 539 595 573
rect 629 539 652 573
rect 583 536 652 539
rect 461 414 535 536
rect 461 380 487 414
rect 521 380 535 414
rect 461 368 535 380
rect 565 368 652 536
rect 682 580 741 592
rect 682 546 695 580
rect 729 546 741 580
rect 682 497 741 546
rect 682 463 695 497
rect 729 463 741 497
rect 682 414 741 463
rect 682 380 695 414
rect 729 380 741 414
rect 682 368 741 380
<< ndiffc >>
rect 39 154 73 188
rect 39 86 73 120
rect 139 88 173 122
rect 239 154 273 188
rect 239 86 273 120
rect 339 156 373 190
rect 339 86 373 120
rect 494 152 528 186
rect 594 161 628 195
rect 608 82 642 116
rect 694 176 728 210
rect 694 86 728 120
<< pdiffc >>
rect 39 546 73 580
rect 39 478 73 512
rect 39 410 73 444
rect 227 546 261 580
rect 227 478 261 512
rect 227 410 261 444
rect 327 539 361 573
rect 595 539 629 573
rect 487 380 521 414
rect 695 546 729 580
rect 695 463 729 497
rect 695 380 729 414
<< poly >>
rect 86 592 116 618
rect 170 592 200 618
rect 284 592 314 618
rect 652 592 682 618
rect 535 536 565 562
rect 86 377 116 392
rect 170 377 200 392
rect 284 377 314 392
rect 83 360 116 377
rect 167 360 203 377
rect 44 344 114 360
rect 44 310 60 344
rect 94 310 114 344
rect 44 276 114 310
rect 44 242 60 276
rect 94 242 114 276
rect 44 226 114 242
rect 167 344 233 360
rect 167 310 183 344
rect 217 310 233 344
rect 167 276 233 310
rect 167 242 183 276
rect 217 242 233 276
rect 281 302 317 377
rect 535 353 565 368
rect 652 353 682 368
rect 532 310 568 353
rect 649 330 685 353
rect 617 314 685 330
rect 395 302 461 310
rect 281 294 461 302
rect 281 260 411 294
rect 445 260 461 294
rect 281 244 461 260
rect 503 294 569 310
rect 503 260 519 294
rect 553 260 569 294
rect 617 280 633 314
rect 667 280 685 314
rect 617 264 685 280
rect 503 244 569 260
rect 167 226 233 242
rect 84 202 114 226
rect 198 202 228 226
rect 287 202 317 244
rect 539 222 569 244
rect 653 222 683 264
rect 539 86 569 112
rect 84 48 114 74
rect 198 48 228 74
rect 287 48 317 74
rect 653 48 683 74
<< polycont >>
rect 60 310 94 344
rect 60 242 94 276
rect 183 310 217 344
rect 183 242 217 276
rect 411 260 445 294
rect 519 260 553 294
rect 633 280 667 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 512 89 546
rect 23 478 39 512
rect 73 478 89 512
rect 23 444 89 478
rect 23 410 39 444
rect 73 410 89 444
rect 23 394 89 410
rect 211 580 277 596
rect 211 546 227 580
rect 261 546 277 580
rect 211 512 277 546
rect 311 573 377 649
rect 311 539 327 573
rect 361 539 377 573
rect 311 532 377 539
rect 579 573 645 649
rect 579 539 595 573
rect 629 539 645 573
rect 579 532 645 539
rect 679 580 751 596
rect 679 546 695 580
rect 729 546 751 580
rect 211 478 227 512
rect 261 498 277 512
rect 261 478 645 498
rect 211 464 645 478
rect 211 444 357 464
rect 211 410 227 444
rect 261 410 357 444
rect 211 394 357 410
rect 25 344 110 360
rect 25 310 60 344
rect 94 310 110 344
rect 25 276 110 310
rect 25 242 60 276
rect 94 242 110 276
rect 25 226 110 242
rect 167 344 263 360
rect 167 310 183 344
rect 217 310 263 344
rect 167 276 263 310
rect 167 242 183 276
rect 217 242 263 276
rect 167 226 263 242
rect 323 206 357 394
rect 395 414 538 430
rect 395 380 487 414
rect 521 380 538 414
rect 395 364 538 380
rect 395 294 461 364
rect 611 330 645 464
rect 679 497 751 546
rect 679 463 695 497
rect 729 463 751 497
rect 679 414 751 463
rect 679 380 695 414
rect 729 380 751 414
rect 679 364 751 380
rect 611 314 683 330
rect 395 260 411 294
rect 445 260 461 294
rect 395 244 461 260
rect 23 188 289 192
rect 23 154 39 188
rect 73 158 239 188
rect 73 154 89 158
rect 23 120 89 154
rect 223 154 239 158
rect 273 154 289 188
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 122 189 124
rect 123 88 139 122
rect 173 88 189 122
rect 123 17 189 88
rect 223 120 289 154
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 190 389 206
rect 323 156 339 190
rect 373 156 389 190
rect 323 120 389 156
rect 427 202 461 244
rect 503 294 569 310
rect 503 260 519 294
rect 553 260 569 294
rect 611 280 633 314
rect 667 280 683 314
rect 611 264 683 280
rect 503 236 569 260
rect 717 226 751 364
rect 678 210 751 226
rect 427 186 544 202
rect 427 152 494 186
rect 528 152 544 186
rect 427 136 544 152
rect 578 195 644 202
rect 578 161 594 195
rect 628 161 644 195
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 578 116 644 161
rect 578 82 608 116
rect 642 82 644 116
rect 578 17 644 82
rect 678 176 694 210
rect 728 176 751 210
rect 678 120 751 176
rect 678 86 694 120
rect 728 86 751 120
rect 678 70 751 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21ba_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3420808
string GDS_START 3413480
<< end >>
