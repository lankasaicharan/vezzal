magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 43 49 570 157
rect 0 0 576 49
<< scnmos >>
rect 126 47 156 131
rect 204 47 234 131
rect 282 47 312 131
rect 385 47 415 131
rect 457 47 487 131
<< scpmoshvt >>
rect 95 416 145 616
rect 201 416 251 616
rect 307 416 357 616
rect 421 416 471 616
<< ndiff >>
rect 69 111 126 131
rect 69 77 81 111
rect 115 77 126 111
rect 69 47 126 77
rect 156 47 204 131
rect 234 47 282 131
rect 312 105 385 131
rect 312 71 323 105
rect 357 71 385 105
rect 312 47 385 71
rect 415 47 457 131
rect 487 110 544 131
rect 487 76 498 110
rect 532 76 544 110
rect 487 47 544 76
<< pdiff >>
rect 38 597 95 616
rect 38 563 50 597
rect 84 563 95 597
rect 38 462 95 563
rect 38 428 50 462
rect 84 428 95 462
rect 38 416 95 428
rect 145 604 201 616
rect 145 570 156 604
rect 190 570 201 604
rect 145 530 201 570
rect 145 496 156 530
rect 190 496 201 530
rect 145 416 201 496
rect 251 597 307 616
rect 251 563 262 597
rect 296 563 307 597
rect 251 462 307 563
rect 251 428 262 462
rect 296 428 307 462
rect 251 416 307 428
rect 357 604 421 616
rect 357 570 368 604
rect 402 570 421 604
rect 357 533 421 570
rect 357 499 368 533
rect 402 499 421 533
rect 357 462 421 499
rect 357 428 368 462
rect 402 428 421 462
rect 357 416 421 428
rect 471 597 528 616
rect 471 563 482 597
rect 516 563 528 597
rect 471 462 528 563
rect 471 428 482 462
rect 516 428 528 462
rect 471 416 528 428
<< ndiffc >>
rect 81 77 115 111
rect 323 71 357 105
rect 498 76 532 110
<< pdiffc >>
rect 50 563 84 597
rect 50 428 84 462
rect 156 570 190 604
rect 156 496 190 530
rect 262 563 296 597
rect 262 428 296 462
rect 368 570 402 604
rect 368 499 402 533
rect 368 428 402 462
rect 482 563 516 597
rect 482 428 516 462
<< poly >>
rect 95 616 145 642
rect 201 616 251 642
rect 307 616 357 642
rect 421 616 471 642
rect 95 305 145 416
rect 201 374 251 416
rect 307 374 357 416
rect 21 289 145 305
rect 21 255 37 289
rect 71 275 145 289
rect 193 358 259 374
rect 193 324 209 358
rect 243 324 259 358
rect 193 290 259 324
rect 71 255 87 275
rect 21 221 87 255
rect 193 256 209 290
rect 243 256 259 290
rect 193 240 259 256
rect 307 358 373 374
rect 307 324 323 358
rect 357 324 373 358
rect 307 290 373 324
rect 307 256 323 290
rect 357 256 373 290
rect 307 240 373 256
rect 421 304 471 416
rect 421 288 487 304
rect 421 254 437 288
rect 471 254 487 288
rect 21 187 37 221
rect 71 192 87 221
rect 71 187 156 192
rect 21 162 156 187
rect 126 131 156 162
rect 204 131 234 240
rect 307 176 337 240
rect 421 220 487 254
rect 421 192 437 220
rect 282 146 337 176
rect 385 186 437 192
rect 471 186 487 220
rect 385 162 487 186
rect 282 131 312 146
rect 385 131 415 162
rect 457 131 487 162
rect 126 21 156 47
rect 204 21 234 47
rect 282 21 312 47
rect 385 21 415 47
rect 457 21 487 47
<< polycont >>
rect 37 255 71 289
rect 209 324 243 358
rect 209 256 243 290
rect 323 324 357 358
rect 323 256 357 290
rect 437 254 471 288
rect 37 187 71 221
rect 437 186 471 220
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 34 597 100 613
rect 34 563 50 597
rect 84 563 100 597
rect 34 462 100 563
rect 140 604 206 649
rect 140 570 156 604
rect 190 570 206 604
rect 140 530 206 570
rect 140 496 156 530
rect 190 496 206 530
rect 140 480 206 496
rect 246 597 312 613
rect 246 563 262 597
rect 296 563 312 597
rect 34 428 50 462
rect 84 444 100 462
rect 246 462 312 563
rect 246 444 262 462
rect 84 428 262 444
rect 296 428 312 462
rect 34 410 312 428
rect 352 604 418 649
rect 352 570 368 604
rect 402 570 418 604
rect 352 533 418 570
rect 352 499 368 533
rect 402 499 418 533
rect 352 462 418 499
rect 352 428 368 462
rect 402 428 418 462
rect 352 412 418 428
rect 466 597 557 613
rect 466 563 482 597
rect 516 563 557 597
rect 466 462 557 563
rect 466 428 482 462
rect 516 428 557 462
rect 466 412 557 428
rect 21 289 87 356
rect 21 255 37 289
rect 71 255 87 289
rect 21 221 87 255
rect 21 187 37 221
rect 71 187 87 221
rect 21 171 87 187
rect 123 204 157 410
rect 193 358 263 374
rect 193 324 209 358
rect 243 324 263 358
rect 193 290 263 324
rect 193 256 209 290
rect 243 256 263 290
rect 193 240 263 256
rect 307 358 373 374
rect 307 324 323 358
rect 357 324 373 358
rect 307 290 373 324
rect 307 256 323 290
rect 357 256 373 290
rect 307 240 373 256
rect 421 288 487 304
rect 421 254 437 288
rect 471 254 487 288
rect 421 220 487 254
rect 421 204 437 220
rect 123 186 437 204
rect 471 186 487 220
rect 123 170 487 186
rect 123 135 157 170
rect 65 111 157 135
rect 523 134 557 412
rect 65 77 81 111
rect 115 77 157 111
rect 65 53 157 77
rect 307 105 373 134
rect 307 71 323 105
rect 357 71 373 105
rect 307 17 373 71
rect 409 110 557 134
rect 409 76 498 110
rect 532 76 557 110
rect 409 53 557 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3_lp
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5075988
string GDS_START 5070402
<< end >>
