magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 931 235 1303 241
rect 377 157 1303 235
rect 21 49 1303 157
rect 0 0 1344 49
<< scnmos >>
rect 100 47 130 131
rect 242 47 272 131
rect 460 125 490 209
rect 568 125 598 209
rect 640 125 670 209
rect 726 125 756 209
rect 820 125 850 209
rect 1010 47 1040 215
rect 1082 47 1112 215
rect 1190 47 1220 215
<< scpmoshvt >>
rect 100 465 130 593
rect 240 465 270 593
rect 467 447 497 575
rect 568 447 598 575
rect 640 447 670 575
rect 748 447 778 531
rect 820 447 850 531
rect 996 367 1026 619
rect 1082 367 1112 619
rect 1190 367 1220 619
<< ndiff >>
rect 47 110 100 131
rect 47 76 55 110
rect 89 76 100 110
rect 47 47 100 76
rect 130 105 242 131
rect 130 71 197 105
rect 231 71 242 105
rect 130 47 242 71
rect 272 110 325 131
rect 272 76 283 110
rect 317 76 325 110
rect 272 47 325 76
rect 403 187 460 209
rect 403 153 411 187
rect 445 153 460 187
rect 403 125 460 153
rect 490 177 568 209
rect 490 143 501 177
rect 535 143 568 177
rect 490 125 568 143
rect 598 125 640 209
rect 670 177 726 209
rect 670 143 681 177
rect 715 143 726 177
rect 670 125 726 143
rect 756 125 820 209
rect 850 174 903 209
rect 850 140 861 174
rect 895 140 903 174
rect 850 125 903 140
rect 957 171 1010 215
rect 957 137 965 171
rect 999 137 1010 171
rect 957 103 1010 137
rect 957 69 965 103
rect 999 69 1010 103
rect 957 47 1010 69
rect 1040 47 1082 215
rect 1112 124 1190 215
rect 1112 90 1134 124
rect 1168 90 1190 124
rect 1112 47 1190 90
rect 1220 203 1277 215
rect 1220 169 1235 203
rect 1269 169 1277 203
rect 1220 101 1277 169
rect 1220 67 1235 101
rect 1269 67 1277 101
rect 1220 47 1277 67
<< pdiff >>
rect 938 607 996 619
rect 47 581 100 593
rect 47 547 55 581
rect 89 547 100 581
rect 47 511 100 547
rect 47 477 55 511
rect 89 477 100 511
rect 47 465 100 477
rect 130 553 240 593
rect 130 519 145 553
rect 179 519 240 553
rect 130 465 240 519
rect 270 511 323 593
rect 270 477 281 511
rect 315 477 323 511
rect 270 465 323 477
rect 387 447 467 575
rect 497 565 568 575
rect 497 531 516 565
rect 550 531 568 565
rect 497 447 568 531
rect 598 447 640 575
rect 670 561 728 575
rect 670 527 684 561
rect 718 531 728 561
rect 938 573 946 607
rect 980 573 996 607
rect 938 539 996 573
rect 938 531 946 539
rect 718 527 748 531
rect 670 493 748 527
rect 670 459 684 493
rect 718 459 748 493
rect 670 447 748 459
rect 778 447 820 531
rect 850 507 946 531
rect 850 473 861 507
rect 895 505 946 507
rect 980 505 996 539
rect 895 473 996 505
rect 850 455 996 473
rect 850 447 946 455
rect 387 429 445 447
rect 387 395 399 429
rect 433 395 445 429
rect 387 385 445 395
rect 938 421 946 447
rect 980 421 996 455
rect 938 367 996 421
rect 1026 599 1082 619
rect 1026 565 1037 599
rect 1071 565 1082 599
rect 1026 510 1082 565
rect 1026 476 1037 510
rect 1071 476 1082 510
rect 1026 367 1082 476
rect 1112 571 1190 619
rect 1112 537 1131 571
rect 1165 537 1190 571
rect 1112 367 1190 537
rect 1220 578 1273 619
rect 1220 544 1231 578
rect 1265 544 1273 578
rect 1220 367 1273 544
<< ndiffc >>
rect 55 76 89 110
rect 197 71 231 105
rect 283 76 317 110
rect 411 153 445 187
rect 501 143 535 177
rect 681 143 715 177
rect 861 140 895 174
rect 965 137 999 171
rect 965 69 999 103
rect 1134 90 1168 124
rect 1235 169 1269 203
rect 1235 67 1269 101
<< pdiffc >>
rect 55 547 89 581
rect 55 477 89 511
rect 145 519 179 553
rect 281 477 315 511
rect 516 531 550 565
rect 684 527 718 561
rect 946 573 980 607
rect 684 459 718 493
rect 861 473 895 507
rect 946 505 980 539
rect 399 395 433 429
rect 946 421 980 455
rect 1037 565 1071 599
rect 1037 476 1071 510
rect 1131 537 1165 571
rect 1231 544 1265 578
<< poly >>
rect 996 619 1026 645
rect 1082 619 1112 645
rect 1190 619 1220 645
rect 100 593 130 619
rect 240 593 270 619
rect 467 575 497 601
rect 568 575 598 601
rect 640 575 670 601
rect 100 287 130 465
rect 240 443 270 465
rect 217 413 270 443
rect 748 531 778 557
rect 820 531 850 557
rect 217 401 247 413
rect 181 385 247 401
rect 467 415 497 447
rect 460 385 497 415
rect 181 351 197 385
rect 231 351 247 385
rect 460 365 490 385
rect 181 335 247 351
rect 100 271 175 287
rect 100 237 125 271
rect 159 237 175 271
rect 100 203 175 237
rect 100 169 125 203
rect 159 169 175 203
rect 100 153 175 169
rect 217 183 247 335
rect 289 349 490 365
rect 289 315 305 349
rect 339 315 490 349
rect 568 337 598 447
rect 640 415 670 447
rect 640 399 706 415
rect 640 365 656 399
rect 690 365 706 399
rect 640 349 706 365
rect 289 281 490 315
rect 289 247 305 281
rect 339 247 490 281
rect 532 321 598 337
rect 532 287 548 321
rect 582 287 598 321
rect 748 307 778 447
rect 532 271 598 287
rect 289 231 490 247
rect 217 153 272 183
rect 100 131 130 153
rect 242 131 272 153
rect 358 51 388 231
rect 460 209 490 231
rect 568 209 598 271
rect 646 277 778 307
rect 820 415 850 447
rect 820 399 886 415
rect 820 365 836 399
rect 870 365 886 399
rect 820 331 886 365
rect 820 297 836 331
rect 870 297 886 331
rect 996 303 1026 367
rect 820 281 886 297
rect 931 287 1026 303
rect 646 261 676 277
rect 640 231 676 261
rect 640 209 670 231
rect 726 209 756 235
rect 820 209 850 281
rect 931 253 947 287
rect 981 267 1026 287
rect 1082 303 1112 367
rect 1190 335 1220 367
rect 1190 319 1256 335
rect 1082 287 1148 303
rect 981 253 1040 267
rect 931 237 1040 253
rect 1010 215 1040 237
rect 1082 253 1098 287
rect 1132 253 1148 287
rect 1082 237 1148 253
rect 1190 285 1206 319
rect 1240 285 1256 319
rect 1190 269 1256 285
rect 1082 215 1112 237
rect 1190 215 1220 269
rect 460 99 490 125
rect 568 99 598 125
rect 640 51 670 125
rect 726 103 756 125
rect 100 21 130 47
rect 242 21 272 47
rect 358 21 670 51
rect 712 87 778 103
rect 820 99 850 125
rect 712 53 728 87
rect 762 53 778 87
rect 712 37 778 53
rect 1010 21 1040 47
rect 1082 21 1112 47
rect 1190 21 1220 47
<< polycont >>
rect 197 351 231 385
rect 125 237 159 271
rect 125 169 159 203
rect 305 315 339 349
rect 656 365 690 399
rect 305 247 339 281
rect 548 287 582 321
rect 836 365 870 399
rect 836 297 870 331
rect 947 253 981 287
rect 1098 253 1132 287
rect 1206 285 1240 319
rect 728 53 762 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 39 581 93 597
rect 39 547 55 581
rect 89 547 93 581
rect 39 511 93 547
rect 39 477 55 511
rect 89 477 93 511
rect 137 553 179 649
rect 137 519 145 553
rect 137 503 179 519
rect 213 563 409 597
rect 39 469 93 477
rect 213 469 247 563
rect 39 435 247 469
rect 281 511 341 527
rect 315 477 341 511
rect 281 461 341 477
rect 375 497 409 563
rect 500 565 566 649
rect 859 607 983 649
rect 500 531 516 565
rect 550 531 566 565
rect 668 561 760 577
rect 668 527 684 561
rect 718 527 760 561
rect 375 463 598 497
rect 39 110 91 435
rect 39 76 55 110
rect 89 76 91 110
rect 39 60 91 76
rect 125 271 163 401
rect 159 237 163 271
rect 125 203 163 237
rect 159 169 163 203
rect 125 75 163 169
rect 197 385 265 401
rect 231 351 265 385
rect 197 160 265 351
rect 299 349 341 461
rect 299 315 305 349
rect 339 315 341 349
rect 299 281 341 315
rect 299 247 305 281
rect 339 247 341 281
rect 299 126 341 247
rect 383 395 399 429
rect 433 395 449 429
rect 383 253 449 395
rect 532 321 598 463
rect 668 493 760 527
rect 668 459 684 493
rect 718 459 760 493
rect 668 449 760 459
rect 859 573 946 607
rect 980 573 983 607
rect 859 539 983 573
rect 859 507 946 539
rect 859 473 861 507
rect 895 505 946 507
rect 980 505 983 539
rect 895 473 983 505
rect 859 457 983 473
rect 532 287 548 321
rect 582 287 598 321
rect 640 399 692 415
rect 640 365 656 399
rect 690 365 692 399
rect 640 253 692 365
rect 383 219 692 253
rect 726 247 760 449
rect 930 455 983 457
rect 930 421 946 455
rect 980 421 983 455
rect 820 399 886 415
rect 930 405 983 421
rect 1017 599 1077 615
rect 1017 565 1037 599
rect 1071 565 1077 599
rect 1017 510 1077 565
rect 1115 571 1181 649
rect 1115 537 1131 571
rect 1165 537 1181 571
rect 1115 528 1181 537
rect 1215 578 1327 594
rect 1215 544 1231 578
rect 1265 544 1327 578
rect 1215 528 1327 544
rect 1017 476 1037 510
rect 1071 494 1077 510
rect 1071 476 1240 494
rect 1017 460 1240 476
rect 820 365 836 399
rect 870 371 886 399
rect 1017 371 1051 460
rect 870 365 1051 371
rect 820 337 1051 365
rect 820 331 886 337
rect 820 297 836 331
rect 870 297 886 331
rect 820 281 886 297
rect 931 287 981 303
rect 931 253 947 287
rect 931 247 981 253
rect 383 187 449 219
rect 383 153 411 187
rect 445 153 449 187
rect 383 137 449 153
rect 485 177 551 185
rect 485 143 501 177
rect 535 143 551 177
rect 197 105 241 121
rect 231 71 241 105
rect 197 17 241 71
rect 275 110 341 126
rect 275 76 283 110
rect 317 76 341 110
rect 275 60 341 76
rect 485 17 551 143
rect 585 99 629 219
rect 726 213 981 247
rect 726 185 760 213
rect 665 177 760 185
rect 665 143 681 177
rect 715 143 760 177
rect 665 133 760 143
rect 845 174 911 179
rect 1015 175 1051 337
rect 845 140 861 174
rect 895 140 911 174
rect 585 87 778 99
rect 585 53 728 87
rect 762 53 778 87
rect 585 51 778 53
rect 845 17 911 140
rect 949 171 1051 175
rect 949 137 965 171
rect 999 137 1051 171
rect 1085 287 1148 426
rect 1085 253 1098 287
rect 1132 253 1148 287
rect 1190 319 1240 460
rect 1190 285 1206 319
rect 1190 269 1240 285
rect 1085 168 1148 253
rect 1274 219 1327 528
rect 1218 203 1327 219
rect 1218 169 1235 203
rect 1269 169 1327 203
rect 949 103 1051 137
rect 949 69 965 103
rect 999 69 1051 103
rect 949 65 1051 69
rect 1118 124 1184 134
rect 1118 90 1134 124
rect 1168 90 1184 124
rect 1118 17 1184 90
rect 1218 101 1327 169
rect 1218 67 1235 101
rect 1269 67 1327 101
rect 1218 51 1327 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtn_1
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2712608
string GDS_START 2701360
<< end >>
