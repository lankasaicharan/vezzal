magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3698 1975
<< nwell >>
rect -38 332 2438 704
rect 193 322 1355 332
rect 1147 305 1355 322
<< pwell >>
rect 199 207 481 248
rect 1996 228 2399 248
rect 199 184 593 207
rect 944 184 2399 228
rect 1 49 2399 184
rect 0 0 2400 49
<< scpmos >>
rect 83 508 119 592
rect 285 358 321 582
rect 375 358 411 582
rect 583 456 619 540
rect 683 456 719 540
rect 767 456 803 540
rect 990 456 1026 540
rect 1080 456 1116 540
rect 1233 341 1269 541
rect 1334 392 1370 592
rect 1488 508 1524 592
rect 1572 508 1608 592
rect 1680 508 1716 592
rect 1882 508 1918 592
rect 2084 368 2120 568
rect 2191 368 2227 592
rect 2281 368 2317 592
<< nmoslvt >>
rect 84 74 114 158
rect 282 74 312 222
rect 368 74 398 222
rect 582 74 612 158
rect 751 74 781 158
rect 829 74 859 158
rect 1027 118 1057 202
rect 1105 118 1135 202
rect 1248 74 1278 202
rect 1326 74 1356 202
rect 1459 118 1489 202
rect 1566 118 1596 202
rect 1680 118 1710 202
rect 1881 118 1911 202
rect 2079 94 2109 222
rect 2195 74 2225 222
rect 2281 74 2311 222
<< ndiff >>
rect 225 198 282 222
rect 225 164 237 198
rect 271 164 282 198
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 133 171 158
rect 114 99 125 133
rect 159 99 171 133
rect 114 74 171 99
rect 225 119 282 164
rect 225 85 237 119
rect 271 85 282 119
rect 225 74 282 85
rect 312 186 368 222
rect 312 152 323 186
rect 357 152 368 186
rect 312 116 368 152
rect 312 82 323 116
rect 357 82 368 116
rect 312 74 368 82
rect 398 210 455 222
rect 398 176 409 210
rect 443 176 455 210
rect 398 120 455 176
rect 398 86 409 120
rect 443 86 455 120
rect 398 74 455 86
rect 509 169 567 181
rect 509 135 521 169
rect 555 158 567 169
rect 2022 210 2079 222
rect 970 177 1027 202
rect 555 135 582 158
rect 509 74 582 135
rect 612 134 751 158
rect 612 100 673 134
rect 707 100 751 134
rect 612 74 751 100
rect 781 74 829 158
rect 859 123 916 158
rect 859 89 870 123
rect 904 89 916 123
rect 970 143 982 177
rect 1016 143 1027 177
rect 970 118 1027 143
rect 1057 118 1105 202
rect 1135 190 1248 202
rect 1135 156 1146 190
rect 1180 156 1248 190
rect 1135 120 1248 156
rect 1135 118 1199 120
rect 859 74 916 89
rect 1187 86 1199 118
rect 1233 86 1248 120
rect 1187 74 1248 86
rect 1278 74 1326 202
rect 1356 174 1459 202
rect 1356 140 1390 174
rect 1424 140 1459 174
rect 1356 118 1459 140
rect 1489 118 1566 202
rect 1596 118 1680 202
rect 1710 164 1881 202
rect 1710 130 1721 164
rect 1755 130 1822 164
rect 1856 130 1881 164
rect 1710 118 1881 130
rect 1911 177 1968 202
rect 1911 143 1922 177
rect 1956 143 1968 177
rect 1911 118 1968 143
rect 2022 176 2034 210
rect 2068 176 2079 210
rect 2022 140 2079 176
rect 1356 74 1406 118
rect 2022 106 2034 140
rect 2068 106 2079 140
rect 2022 94 2079 106
rect 2109 210 2195 222
rect 2109 176 2136 210
rect 2170 176 2195 210
rect 2109 120 2195 176
rect 2109 94 2136 120
rect 2124 86 2136 94
rect 2170 86 2195 120
rect 2124 74 2195 86
rect 2225 210 2281 222
rect 2225 176 2236 210
rect 2270 176 2281 210
rect 2225 120 2281 176
rect 2225 86 2236 120
rect 2270 86 2281 120
rect 2225 74 2281 86
rect 2311 210 2373 222
rect 2311 176 2327 210
rect 2361 176 2373 210
rect 2311 120 2373 176
rect 2311 86 2327 120
rect 2361 86 2373 120
rect 2311 74 2373 86
<< pdiff >>
rect 27 567 83 592
rect 27 533 39 567
rect 73 533 83 567
rect 27 508 83 533
rect 119 568 175 592
rect 119 534 129 568
rect 163 534 175 568
rect 119 508 175 534
rect 229 404 285 582
rect 229 370 241 404
rect 275 370 285 404
rect 229 358 285 370
rect 321 563 375 582
rect 321 529 331 563
rect 365 529 375 563
rect 321 358 375 529
rect 411 550 467 582
rect 411 516 421 550
rect 455 516 467 550
rect 411 358 467 516
rect 1160 582 1218 594
rect 818 566 911 578
rect 818 540 847 566
rect 527 515 583 540
rect 527 481 539 515
rect 573 481 583 515
rect 527 456 583 481
rect 619 515 683 540
rect 619 481 639 515
rect 673 481 683 515
rect 619 456 683 481
rect 719 456 767 540
rect 803 532 847 540
rect 881 540 911 566
rect 1160 548 1172 582
rect 1206 548 1218 582
rect 1160 541 1218 548
rect 1284 541 1334 592
rect 1160 540 1233 541
rect 881 532 990 540
rect 803 456 990 532
rect 1026 521 1080 540
rect 1026 487 1036 521
rect 1070 487 1080 521
rect 1026 456 1080 487
rect 1116 456 1233 540
rect 1183 341 1233 456
rect 1269 392 1334 541
rect 1370 580 1488 592
rect 1370 546 1444 580
rect 1478 546 1488 580
rect 1370 527 1488 546
rect 1370 493 1380 527
rect 1414 508 1488 527
rect 1524 508 1572 592
rect 1608 579 1680 592
rect 1608 545 1636 579
rect 1670 545 1680 579
rect 1608 508 1680 545
rect 1716 567 1772 592
rect 1716 533 1726 567
rect 1760 533 1772 567
rect 1716 508 1772 533
rect 1826 573 1882 592
rect 1826 539 1838 573
rect 1872 539 1882 573
rect 1826 508 1882 539
rect 1918 567 1974 592
rect 2135 580 2191 592
rect 2135 568 2147 580
rect 1918 533 1928 567
rect 1962 533 1974 567
rect 1918 508 1974 533
rect 2028 556 2084 568
rect 2028 522 2040 556
rect 2074 522 2084 556
rect 1414 493 1426 508
rect 1370 445 1426 493
rect 1370 411 1380 445
rect 1414 411 1426 445
rect 1370 392 1426 411
rect 1269 341 1319 392
rect 2028 485 2084 522
rect 2028 451 2040 485
rect 2074 451 2084 485
rect 2028 414 2084 451
rect 2028 380 2040 414
rect 2074 380 2084 414
rect 2028 368 2084 380
rect 2120 546 2147 568
rect 2181 546 2191 580
rect 2120 498 2191 546
rect 2120 464 2147 498
rect 2181 464 2191 498
rect 2120 368 2191 464
rect 2227 580 2281 592
rect 2227 546 2237 580
rect 2271 546 2281 580
rect 2227 497 2281 546
rect 2227 463 2237 497
rect 2271 463 2281 497
rect 2227 414 2281 463
rect 2227 380 2237 414
rect 2271 380 2281 414
rect 2227 368 2281 380
rect 2317 580 2373 592
rect 2317 546 2327 580
rect 2361 546 2373 580
rect 2317 497 2373 546
rect 2317 463 2327 497
rect 2361 463 2373 497
rect 2317 414 2373 463
rect 2317 380 2327 414
rect 2361 380 2373 414
rect 2317 368 2373 380
<< ndiffc >>
rect 237 164 271 198
rect 39 99 73 133
rect 125 99 159 133
rect 237 85 271 119
rect 323 152 357 186
rect 323 82 357 116
rect 409 176 443 210
rect 409 86 443 120
rect 521 135 555 169
rect 673 100 707 134
rect 870 89 904 123
rect 982 143 1016 177
rect 1146 156 1180 190
rect 1199 86 1233 120
rect 1390 140 1424 174
rect 1721 130 1755 164
rect 1822 130 1856 164
rect 1922 143 1956 177
rect 2034 176 2068 210
rect 2034 106 2068 140
rect 2136 176 2170 210
rect 2136 86 2170 120
rect 2236 176 2270 210
rect 2236 86 2270 120
rect 2327 176 2361 210
rect 2327 86 2361 120
<< pdiffc >>
rect 39 533 73 567
rect 129 534 163 568
rect 241 370 275 404
rect 331 529 365 563
rect 421 516 455 550
rect 539 481 573 515
rect 639 481 673 515
rect 847 532 881 566
rect 1172 548 1206 582
rect 1036 487 1070 521
rect 1444 546 1478 580
rect 1380 493 1414 527
rect 1636 545 1670 579
rect 1726 533 1760 567
rect 1838 539 1872 573
rect 1928 533 1962 567
rect 2040 522 2074 556
rect 1380 411 1414 445
rect 2040 451 2074 485
rect 2040 380 2074 414
rect 2147 546 2181 580
rect 2147 464 2181 498
rect 2237 546 2271 580
rect 2237 463 2271 497
rect 2237 380 2271 414
rect 2327 546 2361 580
rect 2327 463 2361 497
rect 2327 380 2361 414
<< poly >>
rect 83 592 119 618
rect 482 615 1370 645
rect 285 582 321 608
rect 375 582 411 608
rect 83 398 119 508
rect 83 382 161 398
rect 83 348 111 382
rect 145 348 161 382
rect 83 314 161 348
rect 83 280 111 314
rect 145 280 161 314
rect 285 310 321 358
rect 375 326 411 358
rect 482 326 512 615
rect 583 540 619 566
rect 683 540 719 615
rect 1334 592 1370 615
rect 1488 592 1524 618
rect 1572 592 1608 618
rect 1680 592 1716 618
rect 1882 592 1918 618
rect 767 540 803 566
rect 990 540 1026 566
rect 1080 540 1116 566
rect 1233 541 1269 567
rect 583 410 619 456
rect 683 430 719 456
rect 767 414 803 456
rect 368 310 512 326
rect 83 246 161 280
rect 83 212 111 246
rect 145 212 161 246
rect 260 294 326 310
rect 260 260 276 294
rect 310 260 326 294
rect 260 244 326 260
rect 368 276 405 310
rect 439 276 512 310
rect 557 394 623 410
rect 557 360 573 394
rect 607 360 623 394
rect 767 398 912 414
rect 767 384 862 398
rect 557 342 623 360
rect 846 364 862 384
rect 896 364 912 398
rect 846 348 912 364
rect 557 326 787 342
rect 557 292 573 326
rect 607 292 737 326
rect 771 292 787 326
rect 557 276 787 292
rect 368 260 512 276
rect 282 222 312 244
rect 368 222 398 260
rect 482 228 512 260
rect 83 196 161 212
rect 84 158 114 196
rect 482 198 612 228
rect 582 158 612 198
rect 751 158 781 276
rect 882 246 912 348
rect 990 310 1026 456
rect 1080 424 1116 456
rect 1080 408 1151 424
rect 1080 374 1101 408
rect 1135 374 1151 408
rect 1080 358 1151 374
rect 990 294 1057 310
rect 990 260 1006 294
rect 1040 260 1057 294
rect 882 230 948 246
rect 990 244 1057 260
rect 882 210 898 230
rect 829 196 898 210
rect 932 196 948 230
rect 1027 202 1057 244
rect 1105 202 1135 358
rect 2084 568 2120 594
rect 2191 592 2227 618
rect 2281 592 2317 618
rect 1488 476 1524 508
rect 1458 460 1524 476
rect 1458 426 1474 460
rect 1508 426 1524 460
rect 1572 426 1608 508
rect 1680 430 1716 508
rect 1882 457 1918 508
rect 1828 441 1918 457
rect 1458 410 1524 426
rect 1566 410 1632 426
rect 1334 362 1370 392
rect 1566 376 1582 410
rect 1616 376 1632 410
rect 1233 309 1269 341
rect 1334 332 1489 362
rect 1183 293 1278 309
rect 1183 259 1199 293
rect 1233 259 1278 293
rect 1183 243 1278 259
rect 1248 202 1278 243
rect 1326 274 1392 290
rect 1326 240 1342 274
rect 1376 240 1392 274
rect 1326 224 1392 240
rect 1326 202 1356 224
rect 1459 202 1489 332
rect 1566 342 1632 376
rect 1566 308 1582 342
rect 1616 308 1632 342
rect 1566 274 1632 308
rect 1566 240 1582 274
rect 1616 240 1632 274
rect 1566 224 1632 240
rect 1680 414 1746 430
rect 1680 380 1696 414
rect 1730 380 1746 414
rect 1680 346 1746 380
rect 1680 312 1696 346
rect 1730 312 1746 346
rect 1828 407 1844 441
rect 1878 407 1918 441
rect 1828 373 1918 407
rect 1828 339 1844 373
rect 1878 353 1918 373
rect 2084 353 2120 368
rect 1878 339 2120 353
rect 1828 323 2120 339
rect 2191 326 2227 368
rect 2281 326 2317 368
rect 1680 296 1746 312
rect 1566 202 1596 224
rect 1680 202 1710 296
rect 1881 202 1911 323
rect 2079 222 2109 323
rect 2162 310 2317 326
rect 2162 276 2178 310
rect 2212 276 2317 310
rect 2162 260 2317 276
rect 2195 222 2225 260
rect 2281 222 2311 260
rect 829 180 948 196
rect 829 158 859 180
rect 1027 92 1057 118
rect 1105 92 1135 118
rect 1459 92 1489 118
rect 1566 92 1596 118
rect 1680 92 1710 118
rect 1881 92 1911 118
rect 84 48 114 74
rect 282 48 312 74
rect 368 48 398 74
rect 582 48 612 74
rect 751 48 781 74
rect 829 48 859 74
rect 1248 48 1278 74
rect 1326 48 1356 74
rect 2079 68 2109 94
rect 2195 48 2225 74
rect 2281 48 2311 74
<< polycont >>
rect 111 348 145 382
rect 111 280 145 314
rect 111 212 145 246
rect 276 260 310 294
rect 405 276 439 310
rect 573 360 607 394
rect 862 364 896 398
rect 573 292 607 326
rect 737 292 771 326
rect 1101 374 1135 408
rect 1006 260 1040 294
rect 898 196 932 230
rect 1474 426 1508 460
rect 1582 376 1616 410
rect 1199 259 1233 293
rect 1342 240 1376 274
rect 1582 308 1616 342
rect 1582 240 1616 274
rect 1696 380 1730 414
rect 1696 312 1730 346
rect 1844 407 1878 441
rect 1844 339 1878 373
rect 2178 276 2212 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 23 567 73 596
rect 23 533 39 567
rect 23 472 73 533
rect 113 568 179 649
rect 113 534 129 568
rect 163 534 179 568
rect 113 506 179 534
rect 315 563 381 649
rect 315 529 331 563
rect 365 529 381 563
rect 315 506 381 529
rect 421 578 759 612
rect 421 550 455 578
rect 421 480 455 516
rect 489 515 589 544
rect 489 481 539 515
rect 573 481 589 515
rect 23 446 359 472
rect 489 452 589 481
rect 623 515 691 544
rect 623 481 639 515
rect 673 481 691 515
rect 623 452 691 481
rect 489 446 523 452
rect 23 438 523 446
rect 23 153 57 438
rect 325 412 523 438
rect 95 382 161 398
rect 95 348 111 382
rect 145 348 161 382
rect 95 314 161 348
rect 95 280 111 314
rect 145 280 161 314
rect 95 246 161 280
rect 95 212 111 246
rect 145 212 161 246
rect 95 196 161 212
rect 195 370 241 404
rect 275 378 291 404
rect 275 370 455 378
rect 195 344 455 370
rect 195 202 229 344
rect 389 310 455 344
rect 263 294 355 310
rect 263 260 276 294
rect 310 260 355 294
rect 389 276 405 310
rect 439 276 455 310
rect 389 260 455 276
rect 263 236 355 260
rect 409 210 443 226
rect 195 198 287 202
rect 195 164 237 198
rect 271 164 287 198
rect 23 133 73 153
rect 23 99 39 133
rect 23 79 73 99
rect 109 133 159 153
rect 109 99 125 133
rect 109 17 159 99
rect 195 119 287 164
rect 195 85 237 119
rect 271 85 287 119
rect 195 70 287 85
rect 323 186 373 202
rect 357 152 373 186
rect 323 116 373 152
rect 357 82 373 116
rect 323 17 373 82
rect 409 120 443 176
rect 489 185 523 412
rect 557 394 623 410
rect 557 360 573 394
rect 607 360 623 394
rect 557 326 623 360
rect 557 292 573 326
rect 607 292 623 326
rect 557 276 623 292
rect 489 169 555 185
rect 489 135 521 169
rect 489 119 555 135
rect 409 85 443 86
rect 589 85 623 276
rect 409 51 623 85
rect 657 242 691 452
rect 725 482 759 578
rect 814 582 848 649
rect 814 566 915 582
rect 814 532 847 566
rect 881 532 915 566
rect 814 516 915 532
rect 949 578 1138 612
rect 949 482 983 578
rect 725 448 983 482
rect 1017 521 1070 544
rect 1017 487 1036 521
rect 1017 464 1070 487
rect 1104 498 1138 578
rect 1172 582 1222 649
rect 1206 548 1222 582
rect 1172 532 1222 548
rect 1364 580 1494 596
rect 1364 546 1444 580
rect 1478 546 1494 580
rect 1620 579 1686 649
rect 1364 527 1586 546
rect 1620 545 1636 579
rect 1670 545 1686 579
rect 1620 544 1686 545
rect 1726 567 1776 596
rect 1104 464 1317 498
rect 725 326 783 448
rect 1017 414 1051 464
rect 846 398 1051 414
rect 846 364 862 398
rect 896 364 1051 398
rect 846 348 1051 364
rect 1085 424 1223 430
rect 1085 408 1183 424
rect 1085 374 1101 408
rect 1135 390 1183 408
rect 1217 390 1223 424
rect 1135 374 1223 390
rect 1085 358 1223 374
rect 725 292 737 326
rect 771 292 783 326
rect 725 276 783 292
rect 817 294 1249 314
rect 817 280 1006 294
rect 817 242 851 280
rect 990 260 1006 280
rect 1040 293 1249 294
rect 1040 260 1199 293
rect 990 259 1199 260
rect 1233 259 1249 293
rect 657 208 851 242
rect 885 230 954 246
rect 990 244 1249 259
rect 1183 243 1249 244
rect 1283 290 1317 464
rect 1364 493 1380 527
rect 1414 510 1586 527
rect 1760 533 1776 567
rect 1726 510 1776 533
rect 1822 573 1888 649
rect 1822 539 1838 573
rect 1872 539 1888 573
rect 1822 532 1888 539
rect 1928 567 1978 596
rect 2131 580 2197 649
rect 1962 533 1978 567
rect 1364 445 1414 493
rect 1552 498 1776 510
rect 1364 411 1380 445
rect 1364 358 1414 411
rect 1458 460 1518 476
rect 1552 464 1894 498
rect 1458 426 1474 460
rect 1508 430 1518 460
rect 1828 441 1894 464
rect 1508 426 1532 430
rect 1458 396 1532 426
rect 1364 324 1464 358
rect 1283 274 1392 290
rect 657 134 723 208
rect 885 196 898 230
rect 932 210 954 230
rect 1283 240 1342 274
rect 1376 240 1392 274
rect 1283 224 1392 240
rect 932 196 1032 210
rect 885 177 1032 196
rect 885 176 982 177
rect 954 143 982 176
rect 1016 143 1032 177
rect 657 100 673 134
rect 707 100 723 134
rect 657 80 723 100
rect 854 123 920 142
rect 854 89 870 123
rect 904 89 920 123
rect 954 114 1032 143
rect 1130 190 1249 206
rect 1130 156 1146 190
rect 1180 156 1249 190
rect 1130 120 1249 156
rect 854 17 920 89
rect 1130 86 1199 120
rect 1233 86 1249 120
rect 1130 17 1249 86
rect 1283 90 1317 224
rect 1430 190 1464 324
rect 1365 174 1464 190
rect 1365 140 1390 174
rect 1424 140 1464 174
rect 1365 124 1464 140
rect 1498 90 1532 396
rect 1566 410 1629 426
rect 1566 376 1582 410
rect 1616 376 1629 410
rect 1566 342 1629 376
rect 1566 308 1582 342
rect 1616 308 1629 342
rect 1566 274 1629 308
rect 1663 424 1746 430
rect 1697 414 1746 424
rect 1663 380 1696 390
rect 1730 380 1746 414
rect 1663 346 1746 380
rect 1663 312 1696 346
rect 1730 312 1746 346
rect 1828 407 1844 441
rect 1878 407 1894 441
rect 1828 373 1894 407
rect 1828 339 1844 373
rect 1878 339 1894 373
rect 1828 323 1894 339
rect 1663 296 1746 312
rect 1566 240 1582 274
rect 1616 248 1629 274
rect 1928 248 1978 533
rect 1616 240 1978 248
rect 1566 214 1978 240
rect 1283 56 1532 90
rect 1705 164 1872 180
rect 1705 130 1721 164
rect 1755 130 1822 164
rect 1856 130 1872 164
rect 1705 17 1872 130
rect 1906 177 1978 214
rect 1906 143 1922 177
rect 1956 143 1978 177
rect 1906 127 1978 143
rect 2018 556 2090 572
rect 2018 522 2040 556
rect 2074 522 2090 556
rect 2018 485 2090 522
rect 2018 451 2040 485
rect 2074 451 2090 485
rect 2131 546 2147 580
rect 2181 546 2197 580
rect 2131 498 2197 546
rect 2131 464 2147 498
rect 2181 464 2197 498
rect 2231 580 2293 596
rect 2231 546 2237 580
rect 2271 546 2293 580
rect 2231 497 2293 546
rect 2018 414 2090 451
rect 2231 463 2237 497
rect 2271 463 2293 497
rect 2231 430 2293 463
rect 2018 380 2040 414
rect 2074 380 2090 414
rect 2018 326 2090 380
rect 2137 414 2293 430
rect 2137 380 2237 414
rect 2271 380 2293 414
rect 2137 364 2293 380
rect 2327 580 2377 649
rect 2361 546 2377 580
rect 2327 497 2377 546
rect 2361 463 2377 497
rect 2327 414 2377 463
rect 2361 380 2377 414
rect 2327 364 2377 380
rect 2018 310 2225 326
rect 2018 276 2178 310
rect 2212 276 2225 310
rect 2018 260 2225 276
rect 2018 210 2084 260
rect 2259 226 2293 364
rect 2018 176 2034 210
rect 2068 176 2084 210
rect 2018 140 2084 176
rect 2018 106 2034 140
rect 2068 106 2084 140
rect 2018 90 2084 106
rect 2120 210 2186 226
rect 2120 176 2136 210
rect 2170 176 2186 210
rect 2120 120 2186 176
rect 2120 86 2136 120
rect 2170 86 2186 120
rect 2120 17 2186 86
rect 2220 210 2293 226
rect 2220 176 2236 210
rect 2270 176 2293 210
rect 2220 120 2293 176
rect 2220 86 2236 120
rect 2270 86 2293 120
rect 2220 70 2293 86
rect 2327 210 2377 226
rect 2361 176 2377 210
rect 2327 120 2377 176
rect 2361 86 2377 120
rect 2327 17 2377 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 1183 390 1217 424
rect 1663 414 1697 424
rect 1663 390 1696 414
rect 1696 390 1697 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 1171 424 1229 430
rect 1171 390 1183 424
rect 1217 421 1229 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 1217 393 1663 421
rect 1217 390 1229 393
rect 1171 384 1229 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfstp_2
flabel comment s 895 272 895 272 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 701 306 701 306 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 1663 390 1697 424 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 218984
string GDS_START 202424
<< end >>
