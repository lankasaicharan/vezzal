magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 48 49 876 241
rect 0 0 960 49
<< scnmos >>
rect 127 47 157 215
rect 213 47 243 215
rect 299 47 329 215
rect 385 47 415 215
rect 509 47 539 215
rect 595 47 625 215
rect 681 47 711 215
rect 767 47 797 215
<< scpmoshvt >>
rect 127 367 157 619
rect 213 367 243 619
rect 299 367 329 619
rect 385 367 415 619
rect 523 367 553 619
rect 609 367 639 619
rect 695 367 725 619
rect 781 367 811 619
<< ndiff >>
rect 74 203 127 215
rect 74 169 82 203
rect 116 169 127 203
rect 74 93 127 169
rect 74 59 82 93
rect 116 59 127 93
rect 74 47 127 59
rect 157 192 213 215
rect 157 158 168 192
rect 202 158 213 192
rect 157 103 213 158
rect 157 69 168 103
rect 202 69 213 103
rect 157 47 213 69
rect 243 132 299 215
rect 243 98 254 132
rect 288 98 299 132
rect 243 47 299 98
rect 329 203 385 215
rect 329 169 340 203
rect 374 169 385 203
rect 329 101 385 169
rect 329 67 340 101
rect 374 67 385 101
rect 329 47 385 67
rect 415 183 509 215
rect 415 149 446 183
rect 480 149 509 183
rect 415 93 509 149
rect 415 59 446 93
rect 480 59 509 93
rect 415 47 509 59
rect 539 185 595 215
rect 539 151 550 185
rect 584 151 595 185
rect 539 101 595 151
rect 539 67 550 101
rect 584 67 595 101
rect 539 47 595 67
rect 625 127 681 215
rect 625 93 636 127
rect 670 93 681 127
rect 625 47 681 93
rect 711 203 767 215
rect 711 169 722 203
rect 756 169 767 203
rect 711 101 767 169
rect 711 67 722 101
rect 756 67 767 101
rect 711 47 767 67
rect 797 167 850 215
rect 797 133 808 167
rect 842 133 850 167
rect 797 93 850 133
rect 797 59 808 93
rect 842 59 850 93
rect 797 47 850 59
<< pdiff >>
rect 74 599 127 619
rect 74 565 82 599
rect 116 565 127 599
rect 74 524 127 565
rect 74 490 82 524
rect 116 490 127 524
rect 74 441 127 490
rect 74 407 82 441
rect 116 407 127 441
rect 74 367 127 407
rect 157 599 213 619
rect 157 565 168 599
rect 202 565 213 599
rect 157 509 213 565
rect 157 475 168 509
rect 202 475 213 509
rect 157 367 213 475
rect 243 569 299 619
rect 243 535 254 569
rect 288 535 299 569
rect 243 367 299 535
rect 329 599 385 619
rect 329 565 340 599
rect 374 565 385 599
rect 329 509 385 565
rect 329 475 340 509
rect 374 475 385 509
rect 329 367 385 475
rect 415 599 523 619
rect 415 565 456 599
rect 490 565 523 599
rect 415 525 523 565
rect 415 491 456 525
rect 490 491 523 525
rect 415 441 523 491
rect 415 407 456 441
rect 490 407 523 441
rect 415 367 523 407
rect 553 531 609 619
rect 553 497 564 531
rect 598 497 609 531
rect 553 457 609 497
rect 553 423 564 457
rect 598 423 609 457
rect 553 367 609 423
rect 639 447 695 619
rect 639 413 650 447
rect 684 413 695 447
rect 639 367 695 413
rect 725 539 781 619
rect 725 505 736 539
rect 770 505 781 539
rect 725 367 781 505
rect 811 599 864 619
rect 811 565 822 599
rect 856 565 864 599
rect 811 525 864 565
rect 811 491 822 525
rect 856 491 864 525
rect 811 367 864 491
<< ndiffc >>
rect 82 169 116 203
rect 82 59 116 93
rect 168 158 202 192
rect 168 69 202 103
rect 254 98 288 132
rect 340 169 374 203
rect 340 67 374 101
rect 446 149 480 183
rect 446 59 480 93
rect 550 151 584 185
rect 550 67 584 101
rect 636 93 670 127
rect 722 169 756 203
rect 722 67 756 101
rect 808 133 842 167
rect 808 59 842 93
<< pdiffc >>
rect 82 565 116 599
rect 82 490 116 524
rect 82 407 116 441
rect 168 565 202 599
rect 168 475 202 509
rect 254 535 288 569
rect 340 565 374 599
rect 340 475 374 509
rect 456 565 490 599
rect 456 491 490 525
rect 456 407 490 441
rect 564 497 598 531
rect 564 423 598 457
rect 650 413 684 447
rect 736 505 770 539
rect 822 565 856 599
rect 822 491 856 525
<< poly >>
rect 127 619 157 645
rect 213 619 243 645
rect 299 619 329 645
rect 385 619 415 645
rect 523 619 553 645
rect 609 619 639 645
rect 695 619 725 645
rect 781 619 811 645
rect 127 335 157 367
rect 44 319 157 335
rect 44 285 60 319
rect 94 285 157 319
rect 44 269 157 285
rect 127 215 157 269
rect 213 303 243 367
rect 299 303 329 367
rect 385 335 415 367
rect 523 335 553 367
rect 213 287 329 303
rect 213 253 240 287
rect 274 253 329 287
rect 371 319 437 335
rect 371 285 387 319
rect 421 285 437 319
rect 371 269 437 285
rect 479 319 553 335
rect 479 285 495 319
rect 529 285 553 319
rect 609 303 639 367
rect 695 303 725 367
rect 781 335 811 367
rect 479 269 553 285
rect 595 287 725 303
rect 213 237 329 253
rect 213 215 243 237
rect 299 215 329 237
rect 385 215 415 269
rect 509 215 539 269
rect 595 253 611 287
rect 645 253 725 287
rect 595 237 725 253
rect 767 319 833 335
rect 767 285 783 319
rect 817 285 833 319
rect 767 269 833 285
rect 595 215 625 237
rect 681 215 711 237
rect 767 215 797 269
rect 127 21 157 47
rect 213 21 243 47
rect 299 21 329 47
rect 385 21 415 47
rect 509 21 539 47
rect 595 21 625 47
rect 681 21 711 47
rect 767 21 797 47
<< polycont >>
rect 60 285 94 319
rect 240 253 274 287
rect 387 285 421 319
rect 495 285 529 319
rect 611 253 645 287
rect 783 285 817 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 66 599 125 615
rect 66 565 82 599
rect 116 565 125 599
rect 66 524 125 565
rect 66 490 82 524
rect 116 490 125 524
rect 66 441 125 490
rect 159 599 204 615
rect 159 565 168 599
rect 202 565 204 599
rect 159 509 204 565
rect 238 569 304 649
rect 238 535 254 569
rect 288 535 304 569
rect 238 527 304 535
rect 338 599 383 615
rect 338 565 340 599
rect 374 565 383 599
rect 159 475 168 509
rect 202 493 204 509
rect 338 509 383 565
rect 338 493 340 509
rect 202 475 340 493
rect 374 475 383 509
rect 159 459 383 475
rect 417 599 872 615
rect 417 565 456 599
rect 490 581 822 599
rect 490 565 506 581
rect 417 525 506 565
rect 820 565 822 581
rect 856 565 872 599
rect 417 491 456 525
rect 490 491 506 525
rect 66 407 82 441
rect 116 425 125 441
rect 417 441 506 491
rect 417 425 456 441
rect 116 407 456 425
rect 490 407 506 441
rect 548 539 786 547
rect 548 531 736 539
rect 548 497 564 531
rect 598 505 736 531
rect 770 505 786 539
rect 598 501 786 505
rect 820 525 872 565
rect 598 497 600 501
rect 548 457 600 497
rect 820 491 822 525
rect 856 491 872 525
rect 820 475 872 491
rect 548 423 564 457
rect 598 423 600 457
rect 548 407 600 423
rect 634 447 700 467
rect 634 413 650 447
rect 684 441 700 447
rect 684 413 943 441
rect 634 407 943 413
rect 66 391 448 407
rect 17 323 437 357
rect 17 319 171 323
rect 17 285 60 319
rect 94 285 171 319
rect 371 319 437 323
rect 17 269 171 285
rect 205 253 240 287
rect 274 253 290 287
rect 371 285 387 319
rect 421 285 437 319
rect 479 339 846 373
rect 479 319 545 339
rect 479 285 495 319
rect 529 285 545 319
rect 693 319 846 339
rect 598 287 659 303
rect 205 242 290 253
rect 598 253 611 287
rect 645 253 659 287
rect 693 285 783 319
rect 817 285 846 319
rect 66 203 125 219
rect 324 217 564 251
rect 598 237 659 253
rect 880 235 943 407
rect 324 208 390 217
rect 66 169 82 203
rect 116 169 125 203
rect 66 93 125 169
rect 66 59 82 93
rect 116 59 125 93
rect 66 17 125 59
rect 159 203 390 208
rect 159 192 340 203
rect 159 158 168 192
rect 202 174 340 192
rect 159 103 202 158
rect 338 169 340 174
rect 374 169 390 203
rect 530 203 564 217
rect 718 203 943 235
rect 530 185 722 203
rect 159 69 168 103
rect 159 53 202 69
rect 238 132 304 140
rect 238 98 254 132
rect 288 98 304 132
rect 238 17 304 98
rect 338 101 390 169
rect 338 67 340 101
rect 374 67 390 101
rect 338 51 390 67
rect 430 149 446 183
rect 480 149 496 183
rect 430 93 496 149
rect 430 59 446 93
rect 480 59 496 93
rect 430 17 496 59
rect 530 151 550 185
rect 584 169 722 185
rect 756 201 943 203
rect 756 169 758 201
rect 584 151 586 169
rect 530 101 586 151
rect 530 67 550 101
rect 584 67 586 101
rect 530 51 586 67
rect 620 127 686 135
rect 620 93 636 127
rect 670 93 686 127
rect 620 17 686 93
rect 720 101 758 169
rect 720 67 722 101
rect 756 67 758 101
rect 720 51 758 67
rect 792 133 808 167
rect 842 133 858 167
rect 792 93 858 133
rect 792 59 808 93
rect 842 59 858 93
rect 792 17 858 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4181650
string GDS_START 4173320
<< end >>
